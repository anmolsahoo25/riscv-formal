// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
 `define BSV_ASSIGNMENT_DELAY
`endif

// Single-Ported BRAM
module BRAM1Load(CLK,
                 EN,
                 WE,
                 ADDR,
                 DI,
                 DO
                 );

   parameter                      FILENAME   = "";
   parameter                      PIPELINED  = 0;
   parameter                      ADDR_WIDTH = 1;
   parameter                      DATA_WIDTH = 1;
   parameter                      MEMSIZE    = 1;
   parameter                      BINARY     = 0;

   input                          CLK;
   input                          EN;
   input                          WE;
   input [ADDR_WIDTH-1:0]         ADDR;
   input [DATA_WIDTH-1:0]         DI;
   output [DATA_WIDTH-1:0]        DO;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           RAM[0:MEMSIZE-1];
   reg [DATA_WIDTH-1:0]           DO_R;
   reg [DATA_WIDTH-1:0]           DO_R2;

   // synopsys translate_off
   initial
   begin : init_block
`ifdef BSV_NO_INITIAL_BLOCKS
`else
      DO_R  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DO_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
`endif // !`ifdef BSV_NO_INITIAL_BLOCKS
   end
   // synopsys translate_on

   initial
   begin : init_rom_block
      if (BINARY)
        $readmemb(FILENAME, RAM, 0, MEMSIZE-1);
      else
        $readmemh(FILENAME, RAM, 0, MEMSIZE-1);
   end

   always @(posedge CLK) begin
      if (EN) begin
         if (WE) begin
            RAM[ADDR] <= `BSV_ASSIGNMENT_DELAY DI;
      //      DO_R <= `BSV_ASSIGNMENT_DELAY DI;
         end
         else begin
            DO_R <= `BSV_ASSIGNMENT_DELAY RAM[ADDR];
         end
      end
      DO_R2 <= `BSV_ASSIGNMENT_DELAY DO_R;
   end

   // Output driver
   assign DO = (PIPELINED) ? DO_R2 : DO_R;

endmodule // BRAM1Load
// Copyright (c) 2018 IIT- Madras
// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.

module bram_1r1w(
             clka,
             ena,
             wea,
             addra,
             dina,
             clkb,
             enb,
             addrb,
             doutb
             );

   parameter                      ADDR_WIDTH = 6;
   parameter                      DATA_WIDTH = 256;
   parameter                      MEMSIZE    = 64;

   input                          clka;
   input                          ena;
   input                          wea;
   input [ADDR_WIDTH-1:0]         addra;
   input [DATA_WIDTH-1:0]         dina;

   input                          clkb;
   input                          enb;
   input [ADDR_WIDTH-1:0]         addrb;
   output [DATA_WIDTH-1:0]        doutb;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           ram[0:MEMSIZE-1] /* synthesis syn_ramstyle="no_rw_check" */ ;
   reg [DATA_WIDTH-1:0]           out_reg;

   // synopsys translate_off
   integer                        i;
   initial
   begin : init_block
      for (i = 0; i < MEMSIZE; i = i + 1) begin
         ram[i] = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      end
      out_reg = { ((DATA_WIDTH+1)/2) { 2'b10 } };
   end
   // synopsys translate_on

   always @(posedge clka) begin
      if (ena) begin
         if (wea) begin
            ram[addra] <= dina;
         end
      end
   end

   always @(posedge clkb) begin
      if (enb) begin
        out_reg <= ram[addrb];
      end
   end

   // Output drivers
   assign doutb =  out_reg;

endmodule // BRAM2
// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//

module bram_1rw(
             clka,
             ena,
             wea,
             addra,
             dina,
             douta
             );

   parameter                      ADDR_WIDTH = 1;
   parameter                      DATA_WIDTH = 1;
   parameter                      MEMSIZE    = 1;

   input                          clka;
   input                          ena;
   input                          wea;
   input [ADDR_WIDTH-1:0]         addra;
   input [DATA_WIDTH-1:0]         dina;
   output [DATA_WIDTH-1:0]        douta;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           ram[0:MEMSIZE-1];
   reg [DATA_WIDTH-1:0]           out_reg;

   // synopsys translate_off
   integer                        i;
   initial
   begin : init_block
      for (i = 0; i < MEMSIZE; i = i + 1) begin
         ram[i] = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      end
      out_reg  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
   end
   // synopsys translate_on

   always @(posedge clka) begin
      if (ena) begin
         if (wea) begin
            ram[addra] <= dina;
         end
         else begin
            out_reg <= ram[addra];
         end
      end
   end

   // Output driver
   assign douta=out_reg;

endmodule
// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
 `define BSV_ASSIGNMENT_DELAY
`endif

// Dual-Ported BRAM (WRITE FIRST) with byte enables and ability to load from a file
module BRAM2BELoad(CLKA,
                   ENA,
                   WEA,
                   ADDRA,
                   DIA,
                   DOA,
                   CLKB,
                   ENB,
                   WEB,
                   ADDRB,
                   DIB,
                   DOB
                  );

   parameter                      FILENAME   = "";
   parameter                      PIPELINED  = 0;
   parameter                      ADDR_WIDTH = 1;
   parameter                      DATA_WIDTH = 1;
   parameter                      CHUNKSIZE  = 1;
   parameter                      WE_WIDTH   = 1;
   parameter                      MEMSIZE    = 1;
   parameter                      BINARY     = 0;

   input                          CLKA;
   input                          ENA;
   input [WE_WIDTH-1:0]           WEA;
   input [ADDR_WIDTH-1:0]         ADDRA;
   input [DATA_WIDTH-1:0]         DIA;
   output [DATA_WIDTH-1:0]        DOA;

   input                          CLKB;
   input                          ENB;
   input [WE_WIDTH-1:0]           WEB;
   input [ADDR_WIDTH-1:0]         ADDRB;
   input [DATA_WIDTH-1:0]         DIB;
   output [DATA_WIDTH-1:0]        DOB;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           RAM[0:MEMSIZE-1] /* synthesis syn_ramstyle="no_rw_check" */ ;
   reg [DATA_WIDTH-1:0]           DOA_R;
   reg [DATA_WIDTH-1:0]           DOA_R2;
   reg [DATA_WIDTH-1:0]           DOB_R;
   reg [DATA_WIDTH-1:0]           DOB_R2;

   // synopsys translate_off
   initial
   begin : init_block
`ifdef BSV_NO_INITIAL_BLOCKS
`else
      DOA_R  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOA_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
`endif // !`ifdef BSV_NO_INITIAL_BLOCKS
   end
   // synopsys translate_on

   initial
   begin : init_rom_block
      if (BINARY)
        $readmemb(FILENAME, RAM, 0, MEMSIZE-1);
      else
        $readmemh(FILENAME, RAM, 0, MEMSIZE-1);
   end
   
   // PORT A

   // iverilog does not support the full verilog-2001 language.  This fixes that for simulation.
`ifdef __ICARUS__
   reg [DATA_WIDTH-1:0]  MASKA, IMASKA;
   reg  [DATA_WIDTH-1:0] DATA_A;
   wire [DATA_WIDTH-1:0] DATA_Awr;

   assign DATA_Awr = RAM[ADDRA];

   always @(WEA or DIA or DATA_Awr) begin : combo1
      integer j;
      MASKA  = 0;
      IMASKA = 0;

      for(j = WE_WIDTH-1; j >= 0; j = j - 1) begin
         if (WEA[j]) MASKA = (MASKA << 8) | { { DATA_WIDTH-CHUNKSIZE { 1'b0 } }, { CHUNKSIZE { 1'b1 } } };
         else        MASKA = (MASKA << 8);
      end
      IMASKA = ~MASKA;

      DATA_A = (DATA_Awr & IMASKA) | (DIA & MASKA);
   end

   always @(posedge CLKA) begin
      if (ENA) begin
         if (WEA) begin
            RAM[ADDRA] <= `BSV_ASSIGNMENT_DELAY DATA_A;
            DOA_R      <= `BSV_ASSIGNMENT_DELAY DATA_A;
         end
         else begin
            DOA_R      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRA];
         end
      end
   end
`else
   generate
      genvar i;
      for(i = 0; i < WE_WIDTH; i = i + 1) begin: porta_we
         always @(posedge CLKA) begin
            if (ENA) begin
               if (WEA[i]) begin
                  RAM[ADDRA][((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE] <= `BSV_ASSIGNMENT_DELAY DIA[((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE];
                  DOA_R[((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY DIA[((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE];
               end
               else begin
                  DOA_R[((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRA][((i+1)*CHUNKSIZE)-1 : i*CHUNKSIZE];
               end
            end
         end
      end
   endgenerate
`endif // !`ifdef __ICARUS__

   // PORT B

   // iverilog does not support the full verilog-2001 language.  This fixes that for simulation.
`ifdef __ICARUS__
   reg [DATA_WIDTH-1:0]  MASKB, IMASKB;
   reg  [DATA_WIDTH-1:0] DATA_B;
   wire [DATA_WIDTH-1:0] DATA_Bwr;

   assign DATA_Bwr = RAM[ADDRB];

   always @(WEB or DIB or DATA_Bwr) begin : combo2
      integer j;
      MASKB  = 0;
      IMASKB = 0;

      for(j = WE_WIDTH-1; j >= 0; j = j - 1) begin
         if (WEB[j]) MASKB = (MASKB << 8) | { { DATA_WIDTH-CHUNKSIZE { 1'b0 } }, { CHUNKSIZE { 1'b1 } } };
         else        MASKB = (MASKB << 8);
      end
      IMASKB = ~MASKB;

      DATA_B = (DATA_Bwr & IMASKB) | (DIB & MASKB);
   end

   always @(posedge CLKB) begin
      if (ENB) begin
         if (WEB) begin
            RAM[ADDRB] <= `BSV_ASSIGNMENT_DELAY DATA_B;
            DOB_R      <= `BSV_ASSIGNMENT_DELAY DATA_B;
         end
         else begin
            DOB_R      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRB];
         end
      end
   end
`else
   generate
      genvar k;
      for(k = 0; k < WE_WIDTH; k = k + 1) begin: portb_we
         always @(posedge CLKB) begin
            if (ENB) begin
               if (WEB[k]) begin
                  RAM[ADDRB][((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE] <= `BSV_ASSIGNMENT_DELAY DIB[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
                  DOB_R[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY DIB[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
               end
               else begin
                  DOB_R[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRB][((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
               end
            end
         end
      end
   endgenerate
`endif // !`ifdef __ICARUS__

   // Output drivers
   always @(posedge CLKA) begin
      DOA_R2 <= `BSV_ASSIGNMENT_DELAY DOA_R;
   end

   always @(posedge CLKB) begin
      DOB_R2 <= `BSV_ASSIGNMENT_DELAY DOB_R;
   end

   assign DOA = (PIPELINED) ? DOA_R2 : DOA_R;
   assign DOB = (PIPELINED) ? DOB_R2 : DOB_R;

endmodule // BRAM2BELoad
// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
 `define BSV_ASSIGNMENT_DELAY
`endif

// Dual-Ported BRAM (WRITE FIRST) with byte enables
module BRAM2BE(CLKA,
               ENA,
               WEA,
               ADDRA,
               DIA,
               DOA,
               CLKB,
               ENB,
               WEB,
               ADDRB,
               DIB,
               DOB
              );

   parameter                      PIPELINED  = 0;
   parameter                      ADDR_WIDTH = 1;
   parameter                      DATA_WIDTH = 1;
   parameter                      CHUNKSIZE  = 1;
   parameter                      WE_WIDTH   = 1;
   parameter                      MEMSIZE    = 1;

   input                          CLKA;
   input                          ENA;
   input [WE_WIDTH-1:0]           WEA;
   input [ADDR_WIDTH-1:0]         ADDRA;
   input [DATA_WIDTH-1:0]         DIA;
   output [DATA_WIDTH-1:0]        DOA;

   input                          CLKB;
   input                          ENB;
   input [WE_WIDTH-1:0]           WEB;
   input [ADDR_WIDTH-1:0]         ADDRB;
   input [DATA_WIDTH-1:0]         DIB;
   output [DATA_WIDTH-1:0]        DOB;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           RAM[0:MEMSIZE-1] /* synthesis syn_ramstyle="no_rw_check" */ ;
   reg [DATA_WIDTH-1:0]           DOA_R;
   reg [DATA_WIDTH-1:0]           DOA_R2;
   reg [DATA_WIDTH-1:0]           DOB_R;
   reg [DATA_WIDTH-1:0]           DOB_R2;

`ifdef BSV_NO_INITIAL_BLOCKS
`else
   // synopsys translate_off
   integer                        i;
   initial
   begin : init_block
      for (i = 0; i < MEMSIZE; i = i + 1) begin
         RAM[i] = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      end
      DOA_R  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOA_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R  = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
   end
   // synopsys translate_on
`endif // !`ifdef BSV_NO_INITIAL_BLOCKS

   // PORT A

   // iverilog does not support the full verilog-2001 language.  This fixes that for simulation.
`ifdef __ICARUS__
   reg [DATA_WIDTH-1:0]  MASKA, IMASKA;
   reg  [DATA_WIDTH-1:0] DATA_A;
   wire [DATA_WIDTH-1:0] DATA_Awr;

   assign DATA_Awr = RAM[ADDRA];

   always @(WEA or DIA or DATA_Awr) begin : combo1
      integer j;
      MASKA  = 0;
      IMASKA = 0;

      for(j = WE_WIDTH-1; j >= 0; j = j - 1) begin
         if (WEA[j]) MASKA = (MASKA << 8) | { { DATA_WIDTH-CHUNKSIZE { 1'b0 } }, { CHUNKSIZE { 1'b1 } } };
         else        MASKA = (MASKA << 8);
      end
      IMASKA = ~MASKA;

      DATA_A = (DATA_Awr & IMASKA) | (DIA & MASKA);
   end

   always @(posedge CLKA) begin
      if (ENA) begin
         if (WEA) begin
            RAM[ADDRA] <= `BSV_ASSIGNMENT_DELAY DATA_A;
            DOA_R      <= `BSV_ASSIGNMENT_DELAY DATA_A;
         end
         else begin
            DOA_R      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRA];
         end
      end
   end
`else
   generate
      genvar j;
      for(j = 0; j < WE_WIDTH; j = j + 1) begin: porta_we
         always @(posedge CLKA) begin
            if (ENA) begin
               if (WEA[j]) begin
                  RAM[ADDRA][((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE] <= `BSV_ASSIGNMENT_DELAY DIA[((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE];
                  DOA_R[((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY DIA[((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE];
               end
               else begin
                  DOA_R[((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRA][((j+1)*CHUNKSIZE)-1 : j*CHUNKSIZE];
               end
            end
         end
      end
   endgenerate
`endif // !`ifdef __ICARUS__


   // PORT B

   // iverilog does not support the full verilog-2001 language.  This fixes that for simulation.
`ifdef __ICARUS__
   reg [DATA_WIDTH-1:0]  MASKB, IMASKB;
   reg  [DATA_WIDTH-1:0] DATA_B;
   wire [DATA_WIDTH-1:0] DATA_Bwr;

   assign DATA_Bwr = RAM[ADDRB];

   always @(WEB or DIB or DATA_Bwr) begin : combo2
      integer j;
      MASKB  = 0;
      IMASKB = 0;

      for(j = WE_WIDTH-1; j >= 0; j = j - 1) begin
         if (WEB[j]) MASKB = (MASKB << 8) | { { DATA_WIDTH-CHUNKSIZE { 1'b0 } }, { CHUNKSIZE { 1'b1 } } };
         else        MASKB = (MASKB << 8);
      end
      IMASKB = ~MASKB;

      DATA_B = (DATA_Bwr & IMASKB) | (DIB & MASKB);
   end

   always @(posedge CLKB) begin
      if (ENB) begin
         if (WEB) begin
            RAM[ADDRB] <= `BSV_ASSIGNMENT_DELAY DATA_B;
            DOB_R      <= `BSV_ASSIGNMENT_DELAY DATA_B;
         end
         else begin
            DOB_R      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRB];
         end
      end
   end
`else
   generate
      genvar k;
      for(k = 0; k < WE_WIDTH; k = k + 1) begin: portb_we
         always @(posedge CLKB) begin
            if (ENB) begin
               if (WEB[k]) begin
                  RAM[ADDRB][((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE] <= `BSV_ASSIGNMENT_DELAY DIB[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
                  DOB_R[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY DIB[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
               end
               else begin
                  DOB_R[((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE]      <= `BSV_ASSIGNMENT_DELAY RAM[ADDRB][((k+1)*CHUNKSIZE)-1 : k*CHUNKSIZE];
               end
            end
         end
      end
   endgenerate
`endif // !`ifdef __ICARUS__


   // Output drivers
   always @(posedge CLKA) begin
      DOA_R2 <= `BSV_ASSIGNMENT_DELAY DOA_R;
   end

   always @(posedge CLKB) begin
      DOB_R2 <= `BSV_ASSIGNMENT_DELAY DOB_R;
   end

   assign DOA = (PIPELINED) ? DOA_R2 : DOA_R;
   assign DOB = (PIPELINED) ? DOB_R2 : DOB_R;

endmodule // BRAM2BE
// Copyright (c) 2000-2011 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
 `define BSV_ASSIGNMENT_DELAY
`endif

// Dual-Ported BRAM (WRITE FIRST)
module BRAM2(CLKA,
             ENA,
             WEA,
             ADDRA,
             DIA,
             DOA,
             CLKB,
             ENB,
             WEB,
             ADDRB,
             DIB,
             DOB
             );

   parameter                      PIPELINED  = 0;
   parameter                      ADDR_WIDTH = 1;
   parameter                      DATA_WIDTH = 1;
   parameter                      MEMSIZE    = 1;

   input                          CLKA;
   input                          ENA;
   input                          WEA;
   input [ADDR_WIDTH-1:0]         ADDRA;
   input [DATA_WIDTH-1:0]         DIA;
   output [DATA_WIDTH-1:0]        DOA;

   input                          CLKB;
   input                          ENB;
   input                          WEB;
   input [ADDR_WIDTH-1:0]         ADDRB;
   input [DATA_WIDTH-1:0]         DIB;
   output [DATA_WIDTH-1:0]        DOB;

   (* RAM_STYLE = "BLOCK" *)
   reg [DATA_WIDTH-1:0]           RAM[0:MEMSIZE-1] /* synthesis syn_ramstyle="no_rw_check" */ ;
   reg [DATA_WIDTH-1:0]           DOA_R;
   reg [DATA_WIDTH-1:0]           DOB_R;
   reg [DATA_WIDTH-1:0]           DOA_R2;
   reg [DATA_WIDTH-1:0]           DOB_R2;

`ifdef BSV_NO_INITIAL_BLOCKS
`else
   // synopsys translate_off
   integer                        i;
   initial
   begin : init_block
      for (i = 0; i < MEMSIZE; i = i + 1) begin
         RAM[i] = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      end
      DOA_R = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOA_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
      DOB_R2 = { ((DATA_WIDTH+1)/2) { 2'b10 } };
   end
   // synopsys translate_on
`endif // !`ifdef BSV_NO_INITIAL_BLOCKS

   always @(posedge CLKA) begin
      if (ENA) begin
         if (WEA) begin
            RAM[ADDRA] <= `BSV_ASSIGNMENT_DELAY DIA;
            DOA_R <= `BSV_ASSIGNMENT_DELAY DIA;
         end
         else begin
            DOA_R <= `BSV_ASSIGNMENT_DELAY RAM[ADDRA];
         end
      end
      DOA_R2 <= `BSV_ASSIGNMENT_DELAY DOA_R;
   end

   always @(posedge CLKB) begin
      if (ENB) begin
         if (WEB) begin
            RAM[ADDRB] <= `BSV_ASSIGNMENT_DELAY DIB;
            DOB_R <= `BSV_ASSIGNMENT_DELAY DIB;
         end
         else begin
            DOB_R <= `BSV_ASSIGNMENT_DELAY RAM[ADDRB];
         end
      end
      DOB_R2 <= `BSV_ASSIGNMENT_DELAY DOB_R;
   end

   // Output drivers
   assign DOA = (PIPELINED) ? DOA_R2 : DOA_R;
   assign DOB = (PIPELINED) ? DOB_R2 : DOB_R;

endmodule // BRAM2

// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif

module ClockInverter(CLK_IN, PREEDGE,  CLK_OUT);

   input     CLK_IN;            // input clock
   output    PREEDGE;           // output signal announcing an upcoming edge
   output    CLK_OUT;           // output clock

   wire      CLK_OUT;
   wire      PREEDGE;
   
   assign    CLK_OUT = ! CLK_IN ;
   assign    PREEDGE = 1 ;
   
endmodule // ClockInverter


// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif


// N -bit counter with load, set and 2 increment
module Counter(CLK,
               RST,
               Q_OUT,
               DATA_A, ADDA,
               DATA_B, ADDB,
               DATA_C, SETC,
               DATA_F, SETF);

   parameter width = 1;
   parameter init = 0;

   input                 CLK;
   input                 RST;
   input [width - 1 : 0] DATA_A;
   input                 ADDA;
   input [width - 1 : 0] DATA_B;
   input                 ADDB;
   input [width - 1 : 0] DATA_C;
   input                 SETC;
   input [width - 1 : 0] DATA_F;
   input                 SETF;

   output [width - 1 : 0] Q_OUT;



   reg [width - 1 : 0]    q_state ;

   assign                 Q_OUT = q_state ;

   always@(posedge CLK `BSV_ARESET_EDGE_META) begin
    if (RST == `BSV_RESET_VALUE)
      q_state  <= `BSV_ASSIGNMENT_DELAY init;
    else
      begin
         if ( SETF )
           q_state <= `BSV_ASSIGNMENT_DELAY DATA_F ;
         else
           q_state <= `BSV_ASSIGNMENT_DELAY (SETC ? DATA_C : q_state ) + (ADDA ? DATA_A : {width {1'b0}}) + (ADDB ? DATA_B : {width {1'b0}} ) ;
      end // else: !if(RST == `BSV_RESET_VALUE)
   end // always@ (posedge CLK)

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin
      q_state = {((width + 1)/2){2'b10}} ;
   end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif


// Depth 1 FIFO data size 0!
module FIFO10(CLK,
              RST,
              ENQ,
              FULL_N,
              DEQ,
              EMPTY_N,
              CLR
              );

   parameter guarded = 1;

   input                  CLK;
   input                  RST;
   input                  ENQ;
   input                  DEQ;
   input                  CLR ;

   output                 FULL_N;
   output                 EMPTY_N;

   reg                    empty_reg ;

   assign                 EMPTY_N = empty_reg ;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        empty_reg = 1'b0;
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


   assign FULL_N = !empty_reg;

   always@(posedge CLK `BSV_ARESET_EDGE_META)
     begin
        if (RST == `BSV_RESET_VALUE)
          begin
             empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
          end // if (RST == `BSV_RESET_VALUE)
        else
           begin
              if (CLR)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end
              else if (ENQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
                end
              else if (DEQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end // if (DEQ)
           end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if (RST == ! `BSV_RESET_VALUE)
           begin
              if ( ! empty_reg && DEQ )
                begin
                   deqerror = 1 ;
                   $display( "Warning: FIFO10: %m -- Dequeuing from empty fifo" ) ;
                end
              if ( ! FULL_N && ENQ && (!DEQ || guarded) )
                begin
                   enqerror =  1 ;
                   $display( "Warning: FIFO10: %m -- Enqueuing to a full fifo" ) ;
                end
           end // if (RST == ! `BSV_RESET_VALUE)
     end
   // synopsys translate_on

endmodule





// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_ARESET_EDGE_HEAD `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_HEAD
`endif

// Depth 1 FIFO
module FIFO1(CLK,
             RST,
             D_IN,
             ENQ,
             FULL_N,
             D_OUT,
             DEQ,
             EMPTY_N,
             CLR
             );

   parameter width = 1;
   parameter guarded = 1;
   input                  CLK;
   input                  RST;
   input [width - 1 : 0]  D_IN;
   input                  ENQ;
   input                  DEQ;
   input                  CLR ;

   output                 FULL_N;
   output [width - 1 : 0] D_OUT;
   output                 EMPTY_N;

   reg [width - 1 : 0]    D_OUT;
   reg                    empty_reg ;


   assign                 EMPTY_N = empty_reg ;


`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        D_OUT   = {((width + 1)/2) {2'b10}} ;
        empty_reg = 1'b0 ;
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


   assign FULL_N = !empty_reg;

   always@(posedge CLK `BSV_ARESET_EDGE_META)
     begin
        if (RST == `BSV_RESET_VALUE)
          begin
             empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
          end // if (RST == `BSV_RESET_VALUE)
        else
           begin
              if (CLR)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end // if (CLR)
              else if (ENQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
                end // if (ENQ)
              else if (DEQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end // if (DEQ)
           end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   always@(posedge CLK `BSV_ARESET_EDGE_HEAD)
     begin
`ifdef BSV_RESET_FIFO_HEAD
        if (RST == `BSV_RESET_VALUE)
          begin
             D_OUT <= `BSV_ASSIGNMENT_DELAY {width {1'b0}} ;
          end
        else
`endif
           begin
              if (ENQ)
                D_OUT     <= `BSV_ASSIGNMENT_DELAY D_IN;
           end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if (RST == ! `BSV_RESET_VALUE)
           begin
              if ( ! empty_reg && DEQ )
                begin
                   deqerror = 1 ;
                   $display( "Warning: FIFO1: %m -- Dequeuing from empty fifo" ) ;
                end
              if ( ! FULL_N && ENQ && (!DEQ || guarded) )
                begin
                   enqerror =  1 ;
                   $display( "Warning: FIFO1: %m -- Enqueuing to a full fifo" ) ;
                end
           end // if (RST == ! `BSV_RESET_VALUE)
     end
   // synopsys translate_on

endmodule


// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif


// Depth 2 FIFO  Data width 0
module FIFO20(CLK,
              RST,
              ENQ,
              FULL_N,
              DEQ,
              EMPTY_N,
              CLR
              );
   parameter guarded = 1;

   input  RST;
   input  CLK;
   input  ENQ;
   input  CLR;
   input  DEQ;

   output FULL_N;
   output EMPTY_N;

   reg    empty_reg;
   reg    full_reg;

   assign FULL_N  = full_reg ;
   assign EMPTY_N = empty_reg ;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        empty_reg = 1'b0 ;
        full_reg  = 1'b1 ;
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

   always@(posedge CLK `BSV_ARESET_EDGE_META)
      begin
         if (RST == `BSV_RESET_VALUE)
           begin
              empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
              full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
           end // if (RST == `BSV_RESET_VALUE)
         else
           begin
              if (CLR)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                   full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
                end
              else if (ENQ && !DEQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
                   full_reg  <= `BSV_ASSIGNMENT_DELAY ! empty_reg;
                end // if (ENQ && !DEQ)
              else if (!ENQ && DEQ)
                begin
                   full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
                   empty_reg <= `BSV_ASSIGNMENT_DELAY ! full_reg;
                end // if (!ENQ && DEQ)
           end // else: !if(RST == `BSV_RESET_VALUE)
      end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if (RST == ! `BSV_RESET_VALUE)
          begin
             if ( ! empty_reg && DEQ )
               begin
                  deqerror = 1 ;
                  $display( "Warning: FIFO20: %m -- Dequeuing from empty fifo" ) ;
               end
             if ( ! full_reg && ENQ && (!DEQ || guarded) )
               begin
                  enqerror =  1 ;
                  $display( "Warning: FIFO20: %m -- Enqueuing to a full fifo" ) ;
               end
          end // if (RST == ! `BSV_RESET_VALUE)
     end
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_ARESET_EDGE_HEAD `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_HEAD
`endif

// Depth 2 FIFO
module FIFO2(CLK,
             RST,
             D_IN,
             ENQ,
             FULL_N,
             D_OUT,
             DEQ,
             EMPTY_N,
             CLR);

   parameter width = 1;
   parameter guarded = 1;

   input     CLK ;
   input     RST ;
   input [width - 1 : 0] D_IN;
   input                 ENQ;
   input                 DEQ;
   input                 CLR ;

   output                FULL_N;
   output                EMPTY_N;
   output [width - 1 : 0] D_OUT;

   reg                    full_reg;
   reg                    empty_reg;
   reg [width - 1 : 0]    data0_reg;
   reg [width - 1 : 0]    data1_reg;

   assign                 FULL_N = full_reg ;
   assign                 EMPTY_N = empty_reg ;
   assign                 D_OUT = data0_reg ;


   // Optimize the loading logic since state encoding is not power of 2!
   wire                   d0di = (ENQ && ! empty_reg ) || ( ENQ && DEQ && full_reg ) ;
   wire                   d0d1 = DEQ && ! full_reg ;
   wire                   d0h = ((! DEQ) && (! ENQ )) || (!DEQ && empty_reg ) || ( ! ENQ &&full_reg) ;
   wire                   d1di = ENQ & empty_reg ;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        data0_reg   = {((width + 1)/2) {2'b10}} ;
        data1_reg  = {((width + 1)/2) {2'b10}} ;
        empty_reg = 1'b0;
        full_reg  = 1'b1;
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

   always@(posedge CLK `BSV_ARESET_EDGE_META)
     begin
        if (RST == `BSV_RESET_VALUE)
          begin
             empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
             full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
          end // if (RST == `BSV_RESET_VALUE)
        else
          begin
             if (CLR)
               begin
                  empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                  full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
               end // if (CLR)
             else if ( ENQ && ! DEQ ) // just enq
               begin
                  empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  full_reg <= `BSV_ASSIGNMENT_DELAY ! empty_reg ;
               end
             else if ( DEQ && ! ENQ )
               begin
                  full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  empty_reg <= `BSV_ASSIGNMENT_DELAY ! full_reg;
               end // if ( DEQ && ! ENQ )
          end // else: !if(RST == `BSV_RESET_VALUE)

     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)


   always@(posedge CLK `BSV_ARESET_EDGE_HEAD)
     begin
`ifdef BSV_RESET_FIFO_HEAD
        if (RST == `BSV_RESET_VALUE)
          begin
             data0_reg <= `BSV_ASSIGNMENT_DELAY {width {1'b0}} ;
             data1_reg <= `BSV_ASSIGNMENT_DELAY {width {1'b0}} ;
          end
        else
`endif
          begin
             data0_reg  <= `BSV_ASSIGNMENT_DELAY
                           {width{d0di}} & D_IN | {width{d0d1}} & data1_reg | {width{d0h}} & data0_reg ;
             data1_reg <= `BSV_ASSIGNMENT_DELAY
                          d1di ? D_IN : data1_reg ;
          end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)



   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if (RST == ! `BSV_RESET_VALUE)
          begin
             if ( ! empty_reg && DEQ )
               begin
                  deqerror =  1;
                  $display( "Warning: FIFO2: %m -- Dequeuing from empty fifo" ) ;
               end
             if ( ! full_reg && ENQ && (!DEQ || guarded) )
               begin
                  enqerror = 1;
                  $display( "Warning: FIFO2: %m -- Enqueuing to a full fifo" ) ;
               end
          end
     end // always@ (posedge CLK)
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_ARESET_EDGE_HEAD `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_HEAD
`endif

// Depth 1 FIFO
// Allows simultaneous ENQ and DEQ (at the expense of potentially
// causing combinational loops).
module FIFOL1(CLK,
              RST,
              D_IN,
              ENQ,
              FULL_N,
              D_OUT,
              DEQ,
              EMPTY_N,
              CLR);

   parameter             width = 1;

   input                 CLK;
   input                 RST;

   input [width - 1 : 0] D_IN;
   input                 ENQ;
   input                 DEQ;
   input                 CLR ;

   output                FULL_N;
   output                 EMPTY_N;
   output [width - 1 : 0] D_OUT;



   reg                    empty_reg ;
   reg [width - 1 : 0]    D_OUT;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        D_OUT     <= `BSV_ASSIGNMENT_DELAY {((width + 1)/2) {2'b10}} ;
        empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


   assign FULL_N = !empty_reg || DEQ;
   assign EMPTY_N = empty_reg ;

   always@(posedge CLK `BSV_ARESET_EDGE_META)
     begin
        if (RST == `BSV_RESET_VALUE)
           begin
             empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
           end
        else
           begin
              if (CLR)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end
              else if (ENQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
                end
              else if (DEQ)
                begin
                   empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
                end // if (DEQ)
           end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   always@(posedge CLK `BSV_ARESET_EDGE_HEAD)
     begin
`ifdef BSV_RESET_FIFO_HEAD
        if (RST == `BSV_RESET_VALUE)
          begin
             D_OUT <= `BSV_ASSIGNMENT_DELAY {width {1'b0}} ;
          end
        else
`endif
          begin
              if (ENQ)
                D_OUT     <= `BSV_ASSIGNMENT_DELAY D_IN;
           end // else: !if(RST == `BSV_RESET_VALUE)
     end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if ( ! empty_reg && DEQ )
          begin
             deqerror = 1 ;
             $display( "Warning: FIFOL1: %m -- Dequeuing from empty fifo" ) ;
          end
        if ( ! FULL_N && ENQ && ! DEQ)
          begin
             enqerror =  1 ;
             $display( "Warning: FIFOL1: %m -- Enqueuing to a full fifo" ) ;
          end
     end
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


// Bluespec primitive module which allows creation of clocks
// with non-constant periods.  The CLK_IN and COND_IN inputs
// are registered and used to compute the CLK_OUT and
// CLK_GATE_OUT outputs.
module MakeClock ( CLK, RST,
                   CLK_IN, CLK_IN_EN,
                   COND_IN, COND_IN_EN,
                   CLK_VAL_OUT, COND_OUT,
                   CLK_OUT, CLK_GATE_OUT );

   parameter initVal = 0;
   parameter initGate = 1;

   input  CLK;
   input  RST;

   input  CLK_IN;
   input  CLK_IN_EN;
   input  COND_IN;
   input  COND_IN_EN;

   output CLK_VAL_OUT;
   output COND_OUT;
   output CLK_OUT;
   output CLK_GATE_OUT;

   reg current_clk;
   reg CLK_VAL_OUT;
   reg current_gate;
   reg new_gate;

   // The use of blocking assignment within this block insures
   // that the clock generated from the generate clock (current_clK) occurs before any
   // LHS of nonblocking assigments also from CLKoccur.
   // Basically, this insures that CLK_OUT and CLK occur within
   // the same phase of the execution cycle,  before any state
   // updates occur. see
   // http://www.sunburst-design.com/papers/CummingsSNUG2002Boston_NBAwithDelays.pdf
   always @(posedge CLK or `BSV_RESET_EDGE RST)
   begin
     if (RST == `BSV_RESET_VALUE)
     begin
       current_clk = initVal;
     end
     else
     begin
       if (CLK_IN_EN)
         current_clk = CLK_IN;
     end
   end

   // Duplicate flop for DRC -- clocks cannot be used as data
   always @(posedge CLK or `BSV_RESET_EDGE RST)
   begin
     if (RST == `BSV_RESET_VALUE)
     begin
       CLK_VAL_OUT <=  `BSV_ASSIGNMENT_DELAY initVal;
     end
     else
     begin
       if (CLK_IN_EN)
         CLK_VAL_OUT <=  `BSV_ASSIGNMENT_DELAY CLK_IN;
     end
   end

   always @(posedge CLK or `BSV_RESET_EDGE RST)
   begin
     if (RST == `BSV_RESET_VALUE)
       new_gate   <=  `BSV_ASSIGNMENT_DELAY initGate;
     else
     begin
       if (COND_IN_EN)
         new_gate <=  `BSV_ASSIGNMENT_DELAY  COND_IN;
     end
   end


   // Use latch to avoid glitches
   // Gate can only change when clock is low
   // There remains a fundamental race condition in this design, which
   // is triggered when the current_clk rises and the the new_gate
   // changes.  We recommend to avoid changing the gate in the same
   // cycle when the clock rises.
   always @( current_clk or new_gate )
     begin
        if (current_clk == 1'b0)
          current_gate  <= `BSV_ASSIGNMENT_DELAY new_gate ;
     end

   assign CLK_OUT      = current_clk && current_gate;
   assign CLK_GATE_OUT = current_gate;
   assign COND_OUT     = new_gate;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin
      #0 ;
      current_clk  = 1'b0 ;
      current_gate = 1'b1 ;
      new_gate     = 1'b1 ;
      CLK_VAL_OUT  = 1'b0;
   end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif



module MakeReset0 (
		  CLK,
		  RST,
                  ASSERT_IN,
		  ASSERT_OUT,

                  OUT_RST
                  );

   parameter          init = 1 ;

   input              CLK ;
   input              RST ;
   input              ASSERT_IN ;
   output             ASSERT_OUT ;

   output             OUT_RST ;

   reg                rst ;

   assign ASSERT_OUT =  rst == `BSV_RESET_VALUE ;

   assign OUT_RST = rst ;

   always@(posedge CLK or `BSV_RESET_EDGE RST) begin
      if (RST == `BSV_RESET_VALUE)
        rst <= `BSV_ASSIGNMENT_DELAY init ? ~ `BSV_RESET_VALUE : `BSV_RESET_VALUE;
      else
        begin
           if (ASSERT_IN)
             rst <= `BSV_ASSIGNMENT_DELAY `BSV_RESET_VALUE;
           else // if (rst == 1'b0)
             rst <= `BSV_ASSIGNMENT_DELAY ~ `BSV_RESET_VALUE;
        end // else: !if(RST == `BSV_RESET_VALUE)
   end // always@ (posedge CLK or `BSV_RESET_EDGE RST)


`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin
      #0 ;
      rst = ~ `BSV_RESET_VALUE ;
   end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule // MakeReset0

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif



module MakeResetA (
		  CLK,
		  RST,
                  ASSERT_IN,
		  ASSERT_OUT,

                  DST_CLK,
                  OUT_RST
                  );

   parameter          RSTDELAY = 2  ; // Width of reset shift reg
   parameter          init = 1 ;

   input              CLK ;
   input              RST ;
   input              ASSERT_IN ;
   output             ASSERT_OUT ;

   input              DST_CLK ;
   output             OUT_RST ;

   reg                rst ;
   wire               OUT_RST ;

   assign ASSERT_OUT =  rst == `BSV_RESET_VALUE ;

   SyncResetA #(RSTDELAY) rstSync (.CLK(DST_CLK),
				   .IN_RST(rst),
				   .OUT_RST(OUT_RST));

   always@(posedge CLK or `BSV_RESET_EDGE RST) begin
      if (RST == `BSV_RESET_VALUE)
        rst <= `BSV_ASSIGNMENT_DELAY init ? ~ `BSV_RESET_VALUE : `BSV_RESET_VALUE ;
      else
        begin
           if (ASSERT_IN)
             rst <= `BSV_ASSIGNMENT_DELAY `BSV_RESET_VALUE;
           else // if (rst == 1'b0)
             rst <= `BSV_ASSIGNMENT_DELAY ~ `BSV_RESET_VALUE;
        end // else: !if(RST == `BSV_RESET_VALUE)
   end // always@ (posedge CLK or `BSV_RESET_EDGE RST)

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin
      #0 ;
      rst = ~ `BSV_RESET_VALUE ;
   end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule // MakeResetA
//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:13 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// inputs                         O   138
// RDY_inputs                     O     1 const
// mv_delayed_output              O    65
// RDY_mv_delayed_output          O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// inputs_fn                      I     4
// inputs_op1                     I    64
// inputs_op2                     I    64
// inputs_op3                     I    64
// inputs_imm_value               I    64
// inputs_inst_type               I     4
// inputs_funct3                  I     3
// inputs_memaccess               I     2
// inputs_word32                  I     1
// inputs_misa_c                  I     1
// inputs_lpc                     I     2
// inputs_tdata1                  I    44
// inputs_tdata2                  I   128
// inputs_tenable                 I     2
// EN_inputs                      I     1
//
// Combinational paths from inputs to outputs:
//   (inputs_fn,
//    inputs_op1,
//    inputs_op2,
//    inputs_op3,
//    inputs_imm_value,
//    inputs_inst_type,
//    inputs_funct3,
//    inputs_memaccess,
//    inputs_word32,
//    inputs_misa_c,
//    inputs_lpc,
//    inputs_tdata1,
//    inputs_tdata2,
//    inputs_tenable,
//    EN_inputs) -> inputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkalu(CLK,
	     RST_N,

	     inputs_fn,
	     inputs_op1,
	     inputs_op2,
	     inputs_op3,
	     inputs_imm_value,
	     inputs_inst_type,
	     inputs_funct3,
	     inputs_memaccess,
	     inputs_word32,
	     inputs_misa_c,
	     inputs_lpc,
	     inputs_tdata1,
	     inputs_tdata2,
	     inputs_tenable,
	     EN_inputs,
	     inputs,
	     RDY_inputs,

	     mv_delayed_output,
	     RDY_mv_delayed_output);
  input  CLK;
  input  RST_N;

  // actionvalue method inputs
  input  [3 : 0] inputs_fn;
  input  [63 : 0] inputs_op1;
  input  [63 : 0] inputs_op2;
  input  [63 : 0] inputs_op3;
  input  [63 : 0] inputs_imm_value;
  input  [3 : 0] inputs_inst_type;
  input  [2 : 0] inputs_funct3;
  input  [1 : 0] inputs_memaccess;
  input  inputs_word32;
  input  inputs_misa_c;
  input  [1 : 0] inputs_lpc;
  input  [43 : 0] inputs_tdata1;
  input  [127 : 0] inputs_tdata2;
  input  [1 : 0] inputs_tenable;
  input  EN_inputs;
  output [137 : 0] inputs;
  output RDY_inputs;

  // value method mv_delayed_output
  output [64 : 0] mv_delayed_output;
  output RDY_mv_delayed_output;

  // signals for module outputs
  wire [137 : 0] inputs;
  wire [64 : 0] mv_delayed_output;
  wire RDY_inputs, RDY_mv_delayed_output;

  // inlined wires
  wire [64 : 0] wr_delayed_output_wget;

  // register rg_wait
  reg rg_wait;
  wire rg_wait_D_IN, rg_wait_EN;

  // ports of submodule muldiv
  wire [137 : 0] muldiv_delayed_output, muldiv_get_inputs;
  wire [63 : 0] muldiv_get_inputs_operand1, muldiv_get_inputs_operand2;
  wire [2 : 0] muldiv_get_inputs_funct3;
  wire muldiv_EN_delayed_output,
       muldiv_EN_get_inputs,
       muldiv_RDY_delayed_output,
       muldiv_get_inputs_word32;

  // rule scheduling signals
  wire CAN_FIRE_RL_capture_delayed_muldivputput,
       CAN_FIRE_inputs,
       WILL_FIRE_RL_capture_delayed_muldivputput,
       WILL_FIRE_inputs;

  // inputs to muxes for submodule ports
  wire MUX_rg_wait_write_1__SEL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d7;
  reg TASK_testplusargs___d8;
  reg TASK_testplusargs___d9;
  reg [63 : 0] v__h355;
  // synopsys translate_on

  // remaining internal signals
  reg [21 : 0] CASE_inputs_tdata1_BITS_21_TO_20_2_inputs_tdat_ETC__q3,
	       CASE_inputs_tdata1_BITS_43_TO_42_2_inputs_tdat_ETC__q2;
  reg [1 : 0] CASE_inputs_memaccess_3_inputs_memaccess_1_inp_ETC__q1;
  wire [137 : 0] fn_alu___d42;

  // actionvalue method inputs
  assign inputs =
	     (inputs_inst_type == 4'd8) ? muldiv_get_inputs : fn_alu___d42 ;
  assign RDY_inputs = 1'd1 ;
  assign CAN_FIRE_inputs = 1'd1 ;
  assign WILL_FIRE_inputs = EN_inputs ;

  // value method mv_delayed_output
  assign mv_delayed_output =
	     { wr_delayed_output_wget[64:1],
	       CAN_FIRE_RL_capture_delayed_muldivputput &&
	       wr_delayed_output_wget[0] } ;
  assign RDY_mv_delayed_output = 1'd1 ;

  // submodule muldiv
  mkmuldiv muldiv(.CLK(CLK),
		  .RST_N(RST_N),
		  .get_inputs_funct3(muldiv_get_inputs_funct3),
		  .get_inputs_operand1(muldiv_get_inputs_operand1),
		  .get_inputs_operand2(muldiv_get_inputs_operand2),
		  .get_inputs_word32(muldiv_get_inputs_word32),
		  .EN_get_inputs(muldiv_EN_get_inputs),
		  .EN_delayed_output(muldiv_EN_delayed_output),
		  .get_inputs(muldiv_get_inputs),
		  .RDY_get_inputs(),
		  .delayed_output(muldiv_delayed_output),
		  .RDY_delayed_output(muldiv_RDY_delayed_output));

  // rule RL_capture_delayed_muldivputput
  assign CAN_FIRE_RL_capture_delayed_muldivputput =
	     muldiv_RDY_delayed_output && rg_wait ;
  assign WILL_FIRE_RL_capture_delayed_muldivputput =
	     CAN_FIRE_RL_capture_delayed_muldivputput ;

  // inputs to muxes for submodule ports
  assign MUX_rg_wait_write_1__SEL_1 =
	     EN_inputs && inputs_inst_type == 4'd8 &&
	     !muldiv_get_inputs[137] ;

  // inlined wires
  assign wr_delayed_output_wget = { muldiv_delayed_output[134:71], 1'd1 } ;

  // register rg_wait
  assign rg_wait_D_IN = MUX_rg_wait_write_1__SEL_1 ;
  assign rg_wait_EN =
	     EN_inputs && inputs_inst_type == 4'd8 &&
	     !muldiv_get_inputs[137] ||
	     WILL_FIRE_RL_capture_delayed_muldivputput ;

  // submodule muldiv
  assign muldiv_get_inputs_funct3 = inputs_funct3 ;
  assign muldiv_get_inputs_operand1 = inputs_op1 ;
  assign muldiv_get_inputs_operand2 = inputs_op2 ;
  assign muldiv_get_inputs_word32 = inputs_word32 ;
  assign muldiv_EN_get_inputs = EN_inputs && inputs_inst_type == 4'd8 ;
  assign muldiv_EN_delayed_output = CAN_FIRE_RL_capture_delayed_muldivputput ;

  // remaining internal signals
  module_fn_alu instance_fn_alu_0(.fn_alu_fn(inputs_fn),
				  .fn_alu_op1(inputs_op1),
				  .fn_alu_op2(inputs_op2),
				  .fn_alu_op3(inputs_op3),
				  .fn_alu_imm_value(inputs_imm_value),
				  .fn_alu_inst_type(inputs_inst_type),
				  .fn_alu_funct3(inputs_funct3),
				  .fn_alu_memaccess(CASE_inputs_memaccess_3_inputs_memaccess_1_inp_ETC__q1),
				  .fn_alu_word32(inputs_word32),
				  .fn_alu_misa_c(inputs_misa_c),
				  .fn_alu_lpc(inputs_lpc),
				  .fn_alu_tdata1({ CASE_inputs_tdata1_BITS_43_TO_42_2_inputs_tdat_ETC__q2,
						   CASE_inputs_tdata1_BITS_21_TO_20_2_inputs_tdat_ETC__q3 }),
				  .fn_alu_tdata2(inputs_tdata2),
				  .fn_alu_tenable(inputs_tenable),
				  .fn_alu(fn_alu___d42));
  always@(inputs_memaccess)
  begin
    case (inputs_memaccess)
      2'd3, 2'd1, 2'd0:
	  CASE_inputs_memaccess_3_inputs_memaccess_1_inp_ETC__q1 =
	      inputs_memaccess;
      default: CASE_inputs_memaccess_3_inputs_memaccess_1_inp_ETC__q1 = 2'd2;
    endcase
  end
  always@(inputs_tdata1)
  begin
    case (inputs_tdata1[43:42])
      2'd2, 2'd1, 2'd0:
	  CASE_inputs_tdata1_BITS_43_TO_42_2_inputs_tdat_ETC__q2 =
	      inputs_tdata1[43:22];
      default: CASE_inputs_tdata1_BITS_43_TO_42_2_inputs_tdat_ETC__q2 =
		   { 2'd3,
		     20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(inputs_tdata1)
  begin
    case (inputs_tdata1[21:20])
      2'd2, 2'd1, 2'd0:
	  CASE_inputs_tdata1_BITS_21_TO_20_2_inputs_tdat_ETC__q3 =
	      inputs_tdata1[21:0];
      default: CASE_inputs_tdata1_BITS_21_TO_20_2_inputs_tdat_ETC__q3 =
		   { 2'd3,
		     20'b10101010101010101010 /* unspecified value */  };
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_wait <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_wait_EN) rg_wait <= `BSV_ASSIGNMENT_DELAY rg_wait_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_wait = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput)
	begin
	  TASK_testplusargs___d7 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput)
	begin
	  TASK_testplusargs___d8 = $test$plusargs("malu");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput)
	begin
	  TASK_testplusargs___d9 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput)
	begin
	  v__h355 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput &&
	  (TASK_testplusargs___d7 ||
	   TASK_testplusargs___d8 && TASK_testplusargs___d9))
	$write("[%10d", v__h355, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput &&
	  (TASK_testplusargs___d7 ||
	   TASK_testplusargs___d8 && TASK_testplusargs___d9))
	$write("ALU: Sending delayed Result:%h",
	       muldiv_delayed_output[134:71]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_capture_delayed_muldivputput &&
	  (TASK_testplusargs___d7 ||
	   TASK_testplusargs___d8 && TASK_testplusargs___d9))
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkalu

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:09 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// read_csr                       O    64
// RDY_read_csr                   O     1 const
// RDY_write_csr                  O     1 const
// upd_on_ret                     O    64
// RDY_upd_on_ret                 O     1 const
// upd_on_trap                    O    64
// RDY_upd_on_trap                O     1 const
// RDY_incr_minstret              O     1 const
// mv_csr_decode                  O   152
// RDY_mv_csr_decode              O     1 const
// mv_csr_misa_c                  O     1 reg
// RDY_mv_csr_misa_c              O     1 const
// mv_curr_priv                   O     2
// RDY_mv_curr_priv               O     1 const
// csr_mstatus                    O    64
// RDY_csr_mstatus                O     1 const
// RDY_clint_msip                 O     1 const
// RDY_clint_mtip                 O     1 const
// RDY_clint_mtime                O     1 const
// RDY_ext_interrupt              O     1 const
// mv_interrupt                   O     1
// mv_pmp_cfg                     O    32 reg
// RDY_mv_pmp_cfg                 O     1 const
// mv_pmp_addr                    O   120 reg
// RDY_mv_pmp_addr                O     1 const
// mv_trigger_data1               O    44
// RDY_mv_trigger_data1           O     1 const
// mv_trigger_data2               O   128 reg
// RDY_mv_trigger_data2           O     1 const
// mv_trigger_enable              O     2
// RDY_mv_trigger_enable          O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// read_csr_addr                  I    12
// write_csr_addr                 I    12
// write_csr_word                 I    64
// write_csr_lpc                  I     2
// upd_on_ret_prv                 I     2
// upd_on_trap_cause              I     6
// upd_on_trap_pc                 I    64
// upd_on_trap_tval               I    64
// clint_msip_intrpt              I     1 reg
// clint_mtip_intrpt              I     1 reg
// clint_mtime_c_mtime            I    64 reg
// ext_interrupt_ex_i             I     1 reg
// EN_write_csr                   I     1
// EN_incr_minstret               I     1
// EN_clint_msip                  I     1
// EN_clint_mtip                  I     1
// EN_clint_mtime                 I     1
// EN_ext_interrupt               I     1
// EN_read_csr                    I     1 unused
// EN_upd_on_ret                  I     1
// EN_upd_on_trap                 I     1
//
// Combinational paths from inputs to outputs:
//   read_csr_addr -> read_csr
//   upd_on_ret_prv -> upd_on_ret
//   upd_on_trap_cause -> upd_on_trap
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkcsrfile(CLK,
		 RST_N,

		 read_csr_addr,
		 EN_read_csr,
		 read_csr,
		 RDY_read_csr,

		 write_csr_addr,
		 write_csr_word,
		 write_csr_lpc,
		 EN_write_csr,
		 RDY_write_csr,

		 upd_on_ret_prv,
		 EN_upd_on_ret,
		 upd_on_ret,
		 RDY_upd_on_ret,

		 upd_on_trap_cause,
		 upd_on_trap_pc,
		 upd_on_trap_tval,
		 EN_upd_on_trap,
		 upd_on_trap,
		 RDY_upd_on_trap,

		 EN_incr_minstret,
		 RDY_incr_minstret,

		 mv_csr_decode,
		 RDY_mv_csr_decode,

		 mv_csr_misa_c,
		 RDY_mv_csr_misa_c,

		 mv_curr_priv,
		 RDY_mv_curr_priv,

		 csr_mstatus,
		 RDY_csr_mstatus,

		 clint_msip_intrpt,
		 EN_clint_msip,
		 RDY_clint_msip,

		 clint_mtip_intrpt,
		 EN_clint_mtip,
		 RDY_clint_mtip,

		 clint_mtime_c_mtime,
		 EN_clint_mtime,
		 RDY_clint_mtime,

		 ext_interrupt_ex_i,
		 EN_ext_interrupt,
		 RDY_ext_interrupt,

		 mv_interrupt,

		 mv_pmp_cfg,
		 RDY_mv_pmp_cfg,

		 mv_pmp_addr,
		 RDY_mv_pmp_addr,

		 mv_trigger_data1,
		 RDY_mv_trigger_data1,

		 mv_trigger_data2,
		 RDY_mv_trigger_data2,

		 mv_trigger_enable,
		 RDY_mv_trigger_enable);
  input  CLK;
  input  RST_N;

  // actionvalue method read_csr
  input  [11 : 0] read_csr_addr;
  input  EN_read_csr;
  output [63 : 0] read_csr;
  output RDY_read_csr;

  // action method write_csr
  input  [11 : 0] write_csr_addr;
  input  [63 : 0] write_csr_word;
  input  [1 : 0] write_csr_lpc;
  input  EN_write_csr;
  output RDY_write_csr;

  // actionvalue method upd_on_ret
  input  [1 : 0] upd_on_ret_prv;
  input  EN_upd_on_ret;
  output [63 : 0] upd_on_ret;
  output RDY_upd_on_ret;

  // actionvalue method upd_on_trap
  input  [5 : 0] upd_on_trap_cause;
  input  [63 : 0] upd_on_trap_pc;
  input  [63 : 0] upd_on_trap_tval;
  input  EN_upd_on_trap;
  output [63 : 0] upd_on_trap;
  output RDY_upd_on_trap;

  // action method incr_minstret
  input  EN_incr_minstret;
  output RDY_incr_minstret;

  // value method mv_csr_decode
  output [151 : 0] mv_csr_decode;
  output RDY_mv_csr_decode;

  // value method mv_csr_misa_c
  output mv_csr_misa_c;
  output RDY_mv_csr_misa_c;

  // value method mv_curr_priv
  output [1 : 0] mv_curr_priv;
  output RDY_mv_curr_priv;

  // value method csr_mstatus
  output [63 : 0] csr_mstatus;
  output RDY_csr_mstatus;

  // action method clint_msip
  input  clint_msip_intrpt;
  input  EN_clint_msip;
  output RDY_clint_msip;

  // action method clint_mtip
  input  clint_mtip_intrpt;
  input  EN_clint_mtip;
  output RDY_clint_mtip;

  // action method clint_mtime
  input  [63 : 0] clint_mtime_c_mtime;
  input  EN_clint_mtime;
  output RDY_clint_mtime;

  // action method ext_interrupt
  input  ext_interrupt_ex_i;
  input  EN_ext_interrupt;
  output RDY_ext_interrupt;

  // value method mv_interrupt
  output mv_interrupt;

  // value method mv_pmp_cfg
  output [31 : 0] mv_pmp_cfg;
  output RDY_mv_pmp_cfg;

  // value method mv_pmp_addr
  output [119 : 0] mv_pmp_addr;
  output RDY_mv_pmp_addr;

  // value method mv_trigger_data1
  output [43 : 0] mv_trigger_data1;
  output RDY_mv_trigger_data1;

  // value method mv_trigger_data2
  output [127 : 0] mv_trigger_data2;
  output RDY_mv_trigger_data2;

  // value method mv_trigger_enable
  output [1 : 0] mv_trigger_enable;
  output RDY_mv_trigger_enable;

  // signals for module outputs
  reg [63 : 0] read_csr;
  wire [151 : 0] mv_csr_decode;
  wire [127 : 0] mv_trigger_data2;
  wire [119 : 0] mv_pmp_addr;
  wire [63 : 0] csr_mstatus, upd_on_ret, upd_on_trap;
  wire [43 : 0] mv_trigger_data1;
  wire [31 : 0] mv_pmp_cfg;
  wire [1 : 0] mv_curr_priv, mv_trigger_enable;
  wire RDY_clint_msip,
       RDY_clint_mtime,
       RDY_clint_mtip,
       RDY_csr_mstatus,
       RDY_ext_interrupt,
       RDY_incr_minstret,
       RDY_mv_csr_decode,
       RDY_mv_csr_misa_c,
       RDY_mv_curr_priv,
       RDY_mv_pmp_addr,
       RDY_mv_pmp_cfg,
       RDY_mv_trigger_data1,
       RDY_mv_trigger_data2,
       RDY_mv_trigger_enable,
       RDY_read_csr,
       RDY_upd_on_ret,
       RDY_upd_on_trap,
       RDY_write_csr,
       mv_csr_misa_c,
       mv_interrupt;

  // register ext_ueip
  reg ext_ueip;
  wire ext_ueip_D_IN, ext_ueip_EN;

  // register fflags
  reg [4 : 0] fflags;
  wire [4 : 0] fflags_D_IN;
  wire fflags_EN;

  // register frm
  reg [2 : 0] frm;
  wire [2 : 0] frm_D_IN;
  wire frm_EN;

  // register fs
  reg [1 : 0] fs;
  wire [1 : 0] fs_D_IN;
  wire fs_EN;

  // register mcycle
  reg [63 : 0] mcycle;
  wire [63 : 0] mcycle_D_IN;
  wire mcycle_EN;

  // register minstret
  reg [63 : 0] minstret;
  wire [63 : 0] minstret_D_IN;
  wire minstret_EN;

  // register misa_a
  reg misa_a;
  wire misa_a_D_IN, misa_a_EN;

  // register misa_c
  reg misa_c;
  wire misa_c_D_IN, misa_c_EN;

  // register misa_i
  reg misa_i;
  wire misa_i_D_IN, misa_i_EN;

  // register misa_m
  reg misa_m;
  wire misa_m_D_IN, misa_m_EN;

  // register misa_n
  reg misa_n;
  wire misa_n_D_IN, misa_n_EN;

  // register misa_u
  reg misa_u;
  wire misa_u_D_IN, misa_u_EN;

  // register rg_clint_mtime
  reg [63 : 0] rg_clint_mtime;
  wire [63 : 0] rg_clint_mtime_D_IN;
  wire rg_clint_mtime_EN;

  // register rg_mcause
  reg [4 : 0] rg_mcause;
  wire [4 : 0] rg_mcause_D_IN;
  wire rg_mcause_EN;

  // register rg_mcounteren
  reg [2 : 0] rg_mcounteren;
  wire [2 : 0] rg_mcounteren_D_IN;
  wire rg_mcounteren_EN;

  // register rg_medeleg_l10
  reg [9 : 0] rg_medeleg_l10;
  wire [9 : 0] rg_medeleg_l10_D_IN;
  wire rg_medeleg_l10_EN;

  // register rg_medeleg_m2
  reg [1 : 0] rg_medeleg_m2;
  wire [1 : 0] rg_medeleg_m2_D_IN;
  wire rg_medeleg_m2_EN;

  // register rg_medeleg_u1
  reg rg_medeleg_u1;
  wire rg_medeleg_u1_D_IN, rg_medeleg_u1_EN;

  // register rg_meie
  reg rg_meie;
  wire rg_meie_D_IN, rg_meie_EN;

  // register rg_meip
  reg rg_meip;
  wire rg_meip_D_IN, rg_meip_EN;

  // register rg_mepc
  reg [62 : 0] rg_mepc;
  wire [62 : 0] rg_mepc_D_IN;
  wire rg_mepc_EN;

  // register rg_mideleg
  reg [11 : 0] rg_mideleg;
  wire [11 : 0] rg_mideleg_D_IN;
  wire rg_mideleg_EN;

  // register rg_mie
  reg rg_mie;
  reg rg_mie_D_IN;
  wire rg_mie_EN;

  // register rg_minterrupt
  reg rg_minterrupt;
  wire rg_minterrupt_D_IN, rg_minterrupt_EN;

  // register rg_mode
  reg [1 : 0] rg_mode;
  wire [1 : 0] rg_mode_D_IN;
  wire rg_mode_EN;

  // register rg_mpie
  reg rg_mpie;
  reg rg_mpie_D_IN;
  wire rg_mpie_EN;

  // register rg_mpp
  reg [1 : 0] rg_mpp;
  reg [1 : 0] rg_mpp_D_IN;
  wire rg_mpp_EN;

  // register rg_mprv
  reg rg_mprv;
  wire rg_mprv_D_IN, rg_mprv_EN;

  // register rg_mscratch
  reg [63 : 0] rg_mscratch;
  wire [63 : 0] rg_mscratch_D_IN;
  wire rg_mscratch_EN;

  // register rg_msie
  reg rg_msie;
  wire rg_msie_D_IN, rg_msie_EN;

  // register rg_msip
  reg rg_msip;
  wire rg_msip_D_IN, rg_msip_EN;

  // register rg_mtie
  reg rg_mtie;
  wire rg_mtie_D_IN, rg_mtie_EN;

  // register rg_mtip
  reg rg_mtip;
  wire rg_mtip_D_IN, rg_mtip_EN;

  // register rg_mtval
  reg [63 : 0] rg_mtval;
  wire [63 : 0] rg_mtval_D_IN;
  wire rg_mtval_EN;

  // register rg_mtvec
  reg [61 : 0] rg_mtvec;
  wire [61 : 0] rg_mtvec_D_IN;
  wire rg_mtvec_EN;

  // register rg_prv
  reg [1 : 0] rg_prv;
  wire [1 : 0] rg_prv_D_IN;
  wire rg_prv_EN;

  // register rg_ucause
  reg [4 : 0] rg_ucause;
  wire [4 : 0] rg_ucause_D_IN;
  wire rg_ucause_EN;

  // register rg_ueie
  reg rg_ueie;
  wire rg_ueie_D_IN, rg_ueie_EN;

  // register rg_uepc
  reg [62 : 0] rg_uepc;
  wire [62 : 0] rg_uepc_D_IN;
  wire rg_uepc_EN;

  // register rg_uie
  reg rg_uie;
  reg rg_uie_D_IN;
  wire rg_uie_EN;

  // register rg_uinterrupt
  reg rg_uinterrupt;
  wire rg_uinterrupt_D_IN, rg_uinterrupt_EN;

  // register rg_umode
  reg [1 : 0] rg_umode;
  wire [1 : 0] rg_umode_D_IN;
  wire rg_umode_EN;

  // register rg_upie
  reg rg_upie;
  reg rg_upie_D_IN;
  wire rg_upie_EN;

  // register rg_uscratch
  reg [63 : 0] rg_uscratch;
  wire [63 : 0] rg_uscratch_D_IN;
  wire rg_uscratch_EN;

  // register rg_usie
  reg rg_usie;
  wire rg_usie_D_IN, rg_usie_EN;

  // register rg_usip
  reg rg_usip;
  wire rg_usip_D_IN, rg_usip_EN;

  // register rg_utie
  reg rg_utie;
  wire rg_utie_D_IN, rg_utie_EN;

  // register rg_utip
  reg rg_utip;
  wire rg_utip_D_IN, rg_utip_EN;

  // register rg_utval
  reg [63 : 0] rg_utval;
  wire [63 : 0] rg_utval_D_IN;
  wire rg_utval_EN;

  // register rg_utvec
  reg [61 : 0] rg_utvec;
  wire [61 : 0] rg_utvec_D_IN;
  wire rg_utvec_EN;

  // register soft_ueip
  reg soft_ueip;
  wire soft_ueip_D_IN, soft_ueip_EN;

  // register trigger_index
  reg trigger_index;
  wire trigger_index_D_IN, trigger_index_EN;

  // register v_pmp_addr_0
  reg [29 : 0] v_pmp_addr_0;
  wire [29 : 0] v_pmp_addr_0_D_IN;
  wire v_pmp_addr_0_EN;

  // register v_pmp_addr_1
  reg [29 : 0] v_pmp_addr_1;
  wire [29 : 0] v_pmp_addr_1_D_IN;
  wire v_pmp_addr_1_EN;

  // register v_pmp_addr_2
  reg [29 : 0] v_pmp_addr_2;
  wire [29 : 0] v_pmp_addr_2_D_IN;
  wire v_pmp_addr_2_EN;

  // register v_pmp_addr_3
  reg [29 : 0] v_pmp_addr_3;
  wire [29 : 0] v_pmp_addr_3_D_IN;
  wire v_pmp_addr_3_EN;

  // register v_pmp_cfg_0
  reg [7 : 0] v_pmp_cfg_0;
  wire [7 : 0] v_pmp_cfg_0_D_IN;
  wire v_pmp_cfg_0_EN;

  // register v_pmp_cfg_1
  reg [7 : 0] v_pmp_cfg_1;
  wire [7 : 0] v_pmp_cfg_1_D_IN;
  wire v_pmp_cfg_1_EN;

  // register v_pmp_cfg_2
  reg [7 : 0] v_pmp_cfg_2;
  wire [7 : 0] v_pmp_cfg_2_D_IN;
  wire v_pmp_cfg_2_EN;

  // register v_pmp_cfg_3
  reg [7 : 0] v_pmp_cfg_3;
  wire [7 : 0] v_pmp_cfg_3_D_IN;
  wire v_pmp_cfg_3_EN;

  // register v_tinfo_0
  reg [63 : 0] v_tinfo_0;
  wire [63 : 0] v_tinfo_0_D_IN;
  wire v_tinfo_0_EN;

  // register v_tinfo_1
  reg [63 : 0] v_tinfo_1;
  wire [63 : 0] v_tinfo_1_D_IN;
  wire v_tinfo_1_EN;

  // register v_trig_tdata1_0
  reg [21 : 0] v_trig_tdata1_0;
  wire [21 : 0] v_trig_tdata1_0_D_IN;
  wire v_trig_tdata1_0_EN;

  // register v_trig_tdata1_1
  reg [21 : 0] v_trig_tdata1_1;
  reg [21 : 0] v_trig_tdata1_1_D_IN;
  wire v_trig_tdata1_1_EN;

  // register v_trig_tdata2_0
  reg [63 : 0] v_trig_tdata2_0;
  wire [63 : 0] v_trig_tdata2_0_D_IN;
  wire v_trig_tdata2_0_EN;

  // register v_trig_tdata2_1
  reg [63 : 0] v_trig_tdata2_1;
  wire [63 : 0] v_trig_tdata2_1_D_IN;
  wire v_trig_tdata2_1_EN;

  // register v_trig_tdata3_0
  reg v_trig_tdata3_0;
  wire v_trig_tdata3_0_D_IN, v_trig_tdata3_0_EN;

  // register v_trig_tdata3_1
  reg v_trig_tdata3_1;
  wire v_trig_tdata3_1_D_IN, v_trig_tdata3_1_EN;

  // rule scheduling signals
  wire CAN_FIRE_RL_increment_cycle_counter,
       CAN_FIRE_clint_msip,
       CAN_FIRE_clint_mtime,
       CAN_FIRE_clint_mtip,
       CAN_FIRE_ext_interrupt,
       CAN_FIRE_incr_minstret,
       CAN_FIRE_read_csr,
       CAN_FIRE_upd_on_ret,
       CAN_FIRE_upd_on_trap,
       CAN_FIRE_write_csr,
       WILL_FIRE_RL_increment_cycle_counter,
       WILL_FIRE_clint_msip,
       WILL_FIRE_clint_mtime,
       WILL_FIRE_clint_mtip,
       WILL_FIRE_ext_interrupt,
       WILL_FIRE_incr_minstret,
       WILL_FIRE_read_csr,
       WILL_FIRE_upd_on_ret,
       WILL_FIRE_upd_on_trap,
       WILL_FIRE_write_csr;

  // inputs to muxes for submodule ports
  wire [63 : 0] MUX_mcycle_write_1__VAL_2, MUX_minstret_write_1__VAL_2;
  wire [1 : 0] MUX_rg_prv_write_1__VAL_1, MUX_rg_prv_write_1__VAL_2;
  wire MUX_mcycle_write_1__SEL_1,
       MUX_minstret_write_1__SEL_1,
       MUX_rg_mcause_write_1__SEL_1,
       MUX_rg_mcause_write_1__SEL_2,
       MUX_rg_mepc_write_1__SEL_1,
       MUX_rg_mie_write_1__SEL_1,
       MUX_rg_mie_write_1__SEL_2,
       MUX_rg_mpp_write_1__SEL_3,
       MUX_rg_mtval_write_1__SEL_1,
       MUX_rg_ucause_write_1__SEL_1,
       MUX_rg_uie_write_1__SEL_2,
       MUX_rg_uie_write_1__SEL_3;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d3;
  reg TASK_testplusargs___d4;
  reg TASK_testplusargs___d5;
  reg [63 : 0] v__h3202;
  reg TASK_testplusargs___d9;
  reg TASK_testplusargs___d10;
  reg TASK_testplusargs___d11;
  reg [63 : 0] v__h3355;
  reg TASK_testplusargs___d333;
  reg TASK_testplusargs___d334;
  reg TASK_testplusargs___d335;
  reg [63 : 0] v__h5566;
  reg TASK_testplusargs___d653;
  reg TASK_testplusargs___d654;
  reg TASK_testplusargs___d655;
  reg [63 : 0] v__h10538;
  reg TASK_testplusargs___d659;
  reg TASK_testplusargs___d660;
  reg TASK_testplusargs___d661;
  reg [63 : 0] v__h10688;
  reg TASK_testplusargs___d675;
  reg TASK_testplusargs___d676;
  reg TASK_testplusargs___d677;
  reg [63 : 0] v__h14354;
  reg TASK_testplusargs___d696;
  reg TASK_testplusargs___d697;
  reg TASK_testplusargs___d698;
  reg [63 : 0] v__h14564;
  reg TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d683;
  reg TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d685;
  reg TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d692;
  reg TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d695;
  // synopsys translate_on

  // remaining internal signals
  reg [63 : 0] data___1__h3415, data___1__h3613;
  reg [21 : 0] CASE_v_trig_tdata1_0_BITS_21_TO_20_0_v_trig_td_ETC__q2,
	       CASE_v_trig_tdata1_1_BITS_21_TO_20_0_v_trig_td_ETC__q1;
  reg [5 : 0] CASE_trigger_index_0_v_trig_tdata1_0_BITS_8_TO_ETC__q11;
  reg [3 : 0] CASE_trigger_index_0_v_trig_tdata1_0_BITS_14_T_ETC__q15,
	      CASE_trigger_index_0_v_trig_tdata1_0_BITS_9_TO_ETC__q18,
	      SEL_ARR_v_trig_tdata1_0_4_BITS_5_TO_2_6_v_trig_ETC___d49;
  reg CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q20,
      CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q21,
      CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q22,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_10_1__ETC__q19,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_15_1__ETC__q16,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_16_1__ETC__q17,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_17_1__ETC__q12,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_18_1__ETC__q13,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_19_1__ETC__q14,
      CASE_trigger_index_0_v_trig_tdata1_0_BIT_2_1_v_ETC__q10,
      CASE_trigger_index_0_v_trig_tdata3_0_1_v_trig__ETC__q7,
      CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q5,
      CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q6,
      CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q3,
      CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q4,
      SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45,
      SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d54;
  wire [63 : 0] IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d117,
		IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d118,
		_theResult_____2__h3288,
		data___1__h3506,
		data___1__h3703,
		data___1__h4095,
		data___1__h4119,
		data___1__h4126,
		data___1__h4131,
		data___1__h4147,
		data___1__h4262,
		data___1__h4273,
		data___1__h4282,
		data___1__h4287,
		data___1__h4391,
		data___1__h4458,
		data___1__h4603,
		data___1__h4620,
		data___1__h4637,
		data___1__h4730,
		data___1__h5125,
		data___1__h5131,
		data___1__h5145,
		data___1__h5155,
		data___1__h5188,
		data___1__h5221,
		data___1__h5230,
		data___1__h5232,
		data___1__h5260,
		mv_csr_decode_csr_mstatus__h15074;
  wire [62 : 0] IF_upd_on_ret_prv_EQ_3_41_THEN_IF_misa_c_83_TH_ETC___d652,
		result__h10268,
		result__h10415;
  wire [61 : 0] IF_rg_mode_77_EQ_1_10_AND_upd_on_trap_cause_BI_ETC___d713,
		IF_rg_umode_75_EQ_1_05_AND_upd_on_trap_cause_B_ETC___d709;
  wire [25 : 0] misa__h262;
  wire [15 : 0] SEL_ARR_v_trig_tdata1_0_4_BITS_9_TO_6_6_v_trig_ETC___d91,
		rg_medeleg_u1_CONCAT_0_CONCAT_rg_medeleg_m2_CO_ETC__q9;
  wire [11 : 0] rg_mideleg_SRL_upd_on_trap_cause_BITS_4_TO_0__q8,
		x__h15117,
		x__h15129,
		x__h15156,
		x__h15339;
  wire [10 : 0] SEL_ARR_v_trig_tdata1_0_4_BITS_14_TO_11_4_v_tr_ETC___d90;
  wire [9 : 0] SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d109;
  wire [8 : 0] rg_ueie_79_AND_misa_n_45_AND_soft_ueip_41_OR_e_ETC___d739;
  wire [7 : 0] x__h4122;
  wire [6 : 0] _0_CONCAT_rg_utie_82_AND_misa_n_45_AND_rg_utip__ETC___d738;
  wire [3 : 0] x__h9596, x__h9759;
  wire [2 : 0] SEL_ARR_v_trig_tdata1_0_4_BIT_17_6_v_trig_tdat_ETC___d88;
  wire [1 : 0] x__h14812;
  wire NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691,
       misa_n_45_AND_rg_ueie_79___d247,
       misa_n_45_AND_rg_usie_85___d249,
       misa_n_45_AND_rg_usip_54___d240,
       misa_n_45_AND_rg_utie_82___d248,
       misa_n_45_AND_rg_utip_49___d239,
       misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238,
       r__h4396,
       rg_medeleg_u1_56_CONCAT_0_CONCAT_rg_medeleg_m2_ETC___d673,
       rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d669,
       rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694,
       write_csr_addr_EQ_0x1_35_AND_NOT_fflags_25_EQ__ETC___d453,
       write_csr_addr_EQ_0x2_41_AND_NOT_frm_24_EQ_wri_ETC___d451,
       write_csr_word_BITS_1_TO_0_52_ULT_2___d353,
       x__h4161,
       x__h4195,
       x__h4223,
       y__h4164;

  // actionvalue method read_csr
  always@(read_csr_addr or
	  data___1__h4391 or
	  data___1__h4131 or
	  data___1__h4126 or
	  data___1__h4119 or
	  data___1__h4287 or
	  data___1__h4282 or
	  rg_uscratch or
	  data___1__h4273 or
	  data___1__h4262 or
	  rg_utval or
	  data___1__h4147 or
	  data___1__h5232 or
	  misa_u or
	  misa_n or
	  misa_m or
	  misa_i or
	  misa_c or
	  misa_a or
	  data___1__h5221 or
	  data___1__h5230 or
	  data___1__h5188 or
	  data___1__h5260 or
	  data___1__h5125 or
	  rg_mscratch or
	  data___1__h5145 or
	  data___1__h5131 or
	  rg_mtval or
	  data___1__h5155 or
	  data___1__h4730 or
	  data___1__h4637 or
	  data___1__h4620 or
	  data___1__h4603 or
	  data___1__h4458 or
	  data___1__h4095 or
	  data___1__h3703 or
	  data___1__h3613 or
	  data___1__h3506 or
	  data___1__h3415 or mcycle or rg_clint_mtime or minstret)
  begin
    case (read_csr_addr)
      12'h0: read_csr = data___1__h4391;
      12'h001: read_csr = data___1__h4131;
      12'h002: read_csr = data___1__h4126;
      12'h003: read_csr = data___1__h4119;
      12'h004: read_csr = data___1__h4287;
      12'h005: read_csr = data___1__h4282;
      12'h040: read_csr = rg_uscratch;
      12'h041: read_csr = data___1__h4273;
      12'h042: read_csr = data___1__h4262;
      12'h043: read_csr = rg_utval;
      12'h044: read_csr = data___1__h4147;
      12'h300: read_csr = data___1__h5232;
      12'h301:
	  read_csr =
	      { 43'h40000000000,
		misa_u,
		6'd16,
		misa_n,
		misa_m,
		3'd0,
		misa_i,
		5'd0,
		misa_c,
		1'd0,
		misa_a };
      12'h302: read_csr = data___1__h5221;
      12'h303: read_csr = data___1__h5230;
      12'h304: read_csr = data___1__h5188;
      12'h305: read_csr = data___1__h5260;
      12'h306: read_csr = data___1__h5125;
      12'h340: read_csr = rg_mscratch;
      12'h341: read_csr = data___1__h5145;
      12'h342: read_csr = data___1__h5131;
      12'h343: read_csr = rg_mtval;
      12'h344: read_csr = data___1__h5155;
      12'h3A0: read_csr = data___1__h4730;
      12'h3A2, 12'h7A8, 12'h800: read_csr = 64'd0;
      12'h3B0: read_csr = data___1__h4637;
      12'h3B1: read_csr = data___1__h4620;
      12'h3B2: read_csr = data___1__h4603;
      12'h3B3: read_csr = data___1__h4458;
      12'h7A0: read_csr = data___1__h4095;
      12'h7A1: read_csr = data___1__h3703;
      12'h7A2: read_csr = data___1__h3613;
      12'h7A3: read_csr = data___1__h3506;
      12'h7A4: read_csr = data___1__h3415;
      12'hB00, 12'hC00: read_csr = mcycle;
      12'hB01, 12'hC01: read_csr = rg_clint_mtime;
      12'hB02, 12'hC02: read_csr = minstret;
      default: read_csr = 64'd0;
    endcase
  end
  assign RDY_read_csr = 1'd1 ;
  assign CAN_FIRE_read_csr = 1'd1 ;
  assign WILL_FIRE_read_csr = EN_read_csr ;

  // action method write_csr
  assign RDY_write_csr = 1'd1 ;
  assign CAN_FIRE_write_csr = 1'd1 ;
  assign WILL_FIRE_write_csr = EN_write_csr ;

  // actionvalue method upd_on_ret
  assign upd_on_ret =
	     { IF_upd_on_ret_prv_EQ_3_41_THEN_IF_misa_c_83_TH_ETC___d652,
	       1'b0 } ;
  assign RDY_upd_on_ret = 1'd1 ;
  assign CAN_FIRE_upd_on_ret = 1'd1 ;
  assign WILL_FIRE_upd_on_ret = EN_upd_on_ret ;

  // actionvalue method upd_on_trap
  assign upd_on_trap =
	     { rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ?
		 IF_rg_umode_75_EQ_1_05_AND_upd_on_trap_cause_B_ETC___d709 :
		 IF_rg_mode_77_EQ_1_10_AND_upd_on_trap_cause_BI_ETC___d713,
	       2'b0 } ;
  assign RDY_upd_on_trap = 1'd1 ;
  assign CAN_FIRE_upd_on_trap = 1'd1 ;
  assign WILL_FIRE_upd_on_trap = EN_upd_on_trap ;

  // action method incr_minstret
  assign RDY_incr_minstret = 1'd1 ;
  assign CAN_FIRE_incr_minstret = 1'd1 ;
  assign WILL_FIRE_incr_minstret = EN_incr_minstret ;

  // value method mv_csr_decode
  assign mv_csr_decode =
	     { x__h14812,
	       rg_meip,
	       2'd0,
	       misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238,
	       rg_mtip,
	       2'd0,
	       misa_n_45_AND_rg_utip_49___d239,
	       rg_msip,
	       2'd0,
	       misa_n_45_AND_rg_usip_54___d240,
	       x__h15117,
	       rg_mideleg,
	       x__h15129,
	       x__h15156,
	       misa__h262,
	       mv_csr_decode_csr_mstatus__h15074 } ;
  assign RDY_mv_csr_decode = 1'd1 ;

  // value method mv_csr_misa_c
  assign mv_csr_misa_c = misa_c ;
  assign RDY_mv_csr_misa_c = 1'd1 ;

  // value method mv_curr_priv
  assign mv_curr_priv = (rg_prv == 2'd3) ? rg_prv : 2'd0 ;
  assign RDY_mv_curr_priv = 1'd1 ;

  // value method csr_mstatus
  assign csr_mstatus =
	     { r__h4396,
	       45'd32768,
	       rg_mprv,
	       2'd0,
	       fs,
	       rg_mpp,
	       3'd0,
	       rg_mpie,
	       2'd0,
	       rg_upie,
	       rg_mie,
	       2'd0,
	       rg_uie } ;
  assign RDY_csr_mstatus = 1'd1 ;

  // action method clint_msip
  assign RDY_clint_msip = 1'd1 ;
  assign CAN_FIRE_clint_msip = 1'd1 ;
  assign WILL_FIRE_clint_msip = EN_clint_msip ;

  // action method clint_mtip
  assign RDY_clint_mtip = 1'd1 ;
  assign CAN_FIRE_clint_mtip = 1'd1 ;
  assign WILL_FIRE_clint_mtip = EN_clint_mtip ;

  // action method clint_mtime
  assign RDY_clint_mtime = 1'd1 ;
  assign CAN_FIRE_clint_mtime = 1'd1 ;
  assign WILL_FIRE_clint_mtime = EN_clint_mtime ;

  // action method ext_interrupt
  assign RDY_ext_interrupt = 1'd1 ;
  assign CAN_FIRE_ext_interrupt = 1'd1 ;
  assign WILL_FIRE_ext_interrupt = EN_ext_interrupt ;

  // value method mv_interrupt
  assign mv_interrupt = x__h15339 != 12'd0 ;

  // value method mv_pmp_cfg
  assign mv_pmp_cfg = { v_pmp_cfg_3, v_pmp_cfg_2, v_pmp_cfg_1, v_pmp_cfg_0 } ;
  assign RDY_mv_pmp_cfg = 1'd1 ;

  // value method mv_pmp_addr
  assign mv_pmp_addr =
	     { v_pmp_addr_3, v_pmp_addr_2, v_pmp_addr_1, v_pmp_addr_0 } ;
  assign RDY_mv_pmp_addr = 1'd1 ;

  // value method mv_trigger_data1
  assign mv_trigger_data1 =
	     { CASE_v_trig_tdata1_1_BITS_21_TO_20_0_v_trig_td_ETC__q1,
	       CASE_v_trig_tdata1_0_BITS_21_TO_20_0_v_trig_td_ETC__q2 } ;
  assign RDY_mv_trigger_data1 = 1'd1 ;

  // value method mv_trigger_data2
  assign mv_trigger_data2 = { v_trig_tdata2_1, v_trig_tdata2_0 } ;
  assign RDY_mv_trigger_data2 = 1'd1 ;

  // value method mv_trigger_enable
  assign mv_trigger_enable =
	     { CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q3 &&
	       rg_prv == 2'd3 ||
	       CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q4 &&
	       rg_prv != 2'd3,
	       CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q5 &&
	       rg_prv == 2'd3 ||
	       CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q6 &&
	       rg_prv != 2'd3 } ;
  assign RDY_mv_trigger_enable = 1'd1 ;

  // rule RL_increment_cycle_counter
  assign CAN_FIRE_RL_increment_cycle_counter = 1'd1 ;
  assign WILL_FIRE_RL_increment_cycle_counter = !EN_write_csr ;

  // inputs to muxes for submodule ports
  assign MUX_mcycle_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'hB00 ;
  assign MUX_minstret_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'hB02 ;
  assign MUX_rg_mcause_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'h342 ;
  assign MUX_rg_mcause_write_1__SEL_2 =
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;
  assign MUX_rg_mepc_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'h341 ;
  assign MUX_rg_mie_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'h300 ;
  assign MUX_rg_mie_write_1__SEL_2 = EN_upd_on_ret && upd_on_ret_prv == 2'd3 ;
  assign MUX_rg_mpp_write_1__SEL_3 =
	     EN_write_csr && write_csr_addr == 12'h300 &&
	     (write_csr_word[12:11] == 2'd3 ||
	      write_csr_word[12:11] == 2'd1 ||
	      misa_u && write_csr_word[12:11] == 2'd0) ;
  assign MUX_rg_mtval_write_1__SEL_1 =
	     EN_write_csr && write_csr_addr == 12'h343 ;
  assign MUX_rg_ucause_write_1__SEL_1 =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ;
  assign MUX_rg_uie_write_1__SEL_2 =
	     EN_write_csr &&
	     (write_csr_addr == 12'h300 || write_csr_addr == 12'h0) ;
  assign MUX_rg_uie_write_1__SEL_3 = EN_upd_on_ret && upd_on_ret_prv != 2'd3 ;
  assign MUX_mcycle_write_1__VAL_2 = mcycle + 64'd1 ;
  assign MUX_minstret_write_1__VAL_2 = minstret + 64'd1 ;
  assign MUX_rg_prv_write_1__VAL_1 =
	     (upd_on_ret_prv == 2'd3) ?
	       ((rg_mpp == 2'd3) ? rg_mpp : 2'd0) :
	       2'd0 ;
  assign MUX_rg_prv_write_1__VAL_2 =
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ?
	       2'd0 :
	       2'd3 ;

  // register ext_ueip
  assign ext_ueip_D_IN = ext_interrupt_ex_i ;
  assign ext_ueip_EN = EN_ext_interrupt && rg_prv != 2'd3 ;

  // register fflags
  assign fflags_D_IN = write_csr_word[4:0] ;
  assign fflags_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h001 || write_csr_addr == 12'h003) ;

  // register frm
  assign frm_D_IN =
	     (write_csr_addr == 12'h002) ?
	       write_csr_word[2:0] :
	       write_csr_word[7:5] ;
  assign frm_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h002 || write_csr_addr == 12'h003) ;

  // register fs
  assign fs_D_IN =
	     (write_csr_addr == 12'h300) ? write_csr_word[14:13] : 2'b11 ;
  assign fs_EN =
	     EN_write_csr && write_csr_addr != 12'h301 &&
	     write_csr_addr != 12'h305 &&
	     (write_csr_addr == 12'h300 ||
	      write_csr_addr != 12'h303 && write_csr_addr != 12'h302 &&
	      write_csr_addr != 12'h304 &&
	      write_csr_addr != 12'h344 &&
	      write_csr_addr != 12'hB00 &&
	      write_csr_addr != 12'hB02 &&
	      write_csr_addr != 12'h341 &&
	      write_csr_addr != 12'h343 &&
	      write_csr_addr != 12'h340 &&
	      write_csr_addr != 12'h342 &&
	      write_csr_addr != 12'h306 &&
	      write_csr_addr != 12'h0 &&
	      write_csr_addr != 12'h3A0 &&
	      write_csr_addr != 12'h3A2 &&
	      write_csr_addr != 12'h3B0 &&
	      write_csr_addr != 12'h3B1 &&
	      write_csr_addr != 12'h3B2 &&
	      write_csr_addr != 12'h3B3 &&
	      write_csr_addr != 12'h3B4 &&
	      write_csr_addr != 12'h3B5 &&
	      write_csr_addr != 12'h3B6 &&
	      write_csr_addr != 12'h3B7 &&
	      write_csr_addr != 12'h3B8 &&
	      write_csr_addr != 12'h3B9 &&
	      write_csr_addr != 12'h3BA &&
	      write_csr_addr != 12'h3BB &&
	      write_csr_addr != 12'h3BC &&
	      write_csr_addr != 12'h3BD &&
	      write_csr_addr != 12'h3BE &&
	      write_csr_addr != 12'h3BF &&
	      write_csr_addr != 12'h040 &&
	      write_csr_addr_EQ_0x1_35_AND_NOT_fflags_25_EQ__ETC___d453) ;

  // register mcycle
  assign mcycle_D_IN =
	     MUX_mcycle_write_1__SEL_1 ?
	       write_csr_word :
	       MUX_mcycle_write_1__VAL_2 ;
  assign mcycle_EN =
	     EN_write_csr && write_csr_addr == 12'hB00 ||
	     WILL_FIRE_RL_increment_cycle_counter ;

  // register minstret
  assign minstret_D_IN =
	     MUX_minstret_write_1__SEL_1 ?
	       write_csr_word :
	       MUX_minstret_write_1__VAL_2 ;
  assign minstret_EN =
	     EN_write_csr && write_csr_addr == 12'hB02 || EN_incr_minstret ;

  // register misa_a
  assign misa_a_D_IN = write_csr_word[0] ;
  assign misa_a_EN = EN_write_csr && write_csr_addr == 12'h301 ;

  // register misa_c
  assign misa_c_D_IN = write_csr_word[2] ;
  assign misa_c_EN =
	     EN_write_csr && write_csr_addr == 12'h301 &&
	     (write_csr_word[2] || write_csr_lpc == 2'd0) ;

  // register misa_i
  assign misa_i_D_IN = write_csr_word[8] ;
  assign misa_i_EN = EN_write_csr && write_csr_addr == 12'h301 ;

  // register misa_m
  assign misa_m_D_IN = write_csr_word[12] ;
  assign misa_m_EN = EN_write_csr && write_csr_addr == 12'h301 ;

  // register misa_n
  assign misa_n_D_IN = write_csr_word[13] ;
  assign misa_n_EN = EN_write_csr && write_csr_addr == 12'h301 ;

  // register misa_u
  assign misa_u_D_IN = write_csr_word[20] ;
  assign misa_u_EN = EN_write_csr && write_csr_addr == 12'h301 ;

  // register rg_clint_mtime
  assign rg_clint_mtime_D_IN = clint_mtime_c_mtime ;
  assign rg_clint_mtime_EN = EN_clint_mtime ;

  // register rg_mcause
  assign rg_mcause_D_IN =
	     MUX_rg_mcause_write_1__SEL_1 ?
	       write_csr_word[4:0] :
	       upd_on_trap_cause[4:0] ;
  assign rg_mcause_EN =
	     EN_write_csr && write_csr_addr == 12'h342 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_mcounteren
  assign rg_mcounteren_D_IN = write_csr_word[2:0] ;
  assign rg_mcounteren_EN = EN_write_csr && write_csr_addr == 12'h306 ;

  // register rg_medeleg_l10
  assign rg_medeleg_l10_D_IN = write_csr_word[9:0] ;
  assign rg_medeleg_l10_EN = EN_write_csr && write_csr_addr == 12'h302 ;

  // register rg_medeleg_m2
  assign rg_medeleg_m2_D_IN = write_csr_word[13:12] ;
  assign rg_medeleg_m2_EN = EN_write_csr && write_csr_addr == 12'h302 ;

  // register rg_medeleg_u1
  assign rg_medeleg_u1_D_IN = write_csr_word[15] ;
  assign rg_medeleg_u1_EN = EN_write_csr && write_csr_addr == 12'h302 ;

  // register rg_meie
  assign rg_meie_D_IN = write_csr_word[11] ;
  assign rg_meie_EN = EN_write_csr && write_csr_addr == 12'h304 ;

  // register rg_meip
  assign rg_meip_D_IN = ext_interrupt_ex_i ;
  assign rg_meip_EN = EN_ext_interrupt && rg_prv == 2'd3 ;

  // register rg_mepc
  assign rg_mepc_D_IN =
	     MUX_rg_mepc_write_1__SEL_1 ?
	       write_csr_word[63:1] :
	       upd_on_trap_pc[63:1] ;
  assign rg_mepc_EN =
	     EN_write_csr && write_csr_addr == 12'h341 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_mideleg
  assign rg_mideleg_D_IN = write_csr_word[11:0] ;
  assign rg_mideleg_EN = EN_write_csr && write_csr_addr == 12'h303 ;

  // register rg_mie
  always@(MUX_rg_mie_write_1__SEL_1 or
	  write_csr_word or
	  MUX_rg_mie_write_1__SEL_2 or
	  rg_mpie or MUX_rg_mcause_write_1__SEL_2)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_rg_mie_write_1__SEL_1: rg_mie_D_IN = write_csr_word[3];
      MUX_rg_mie_write_1__SEL_2: rg_mie_D_IN = rg_mpie;
      MUX_rg_mcause_write_1__SEL_2: rg_mie_D_IN = 1'd0;
      default: rg_mie_D_IN = 1'b0 /* unspecified value */ ;
    endcase
  end
  assign rg_mie_EN =
	     EN_write_csr && write_csr_addr == 12'h300 ||
	     EN_upd_on_ret && upd_on_ret_prv == 2'd3 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_minterrupt
  assign rg_minterrupt_D_IN =
	     MUX_rg_mcause_write_1__SEL_1 ?
	       write_csr_word[63] :
	       upd_on_trap_cause[5] ;
  assign rg_minterrupt_EN =
	     EN_write_csr && write_csr_addr == 12'h342 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_mode
  assign rg_mode_D_IN = write_csr_word[1:0] ;
  assign rg_mode_EN =
	     EN_write_csr && write_csr_addr == 12'h305 &&
	     write_csr_word_BITS_1_TO_0_52_ULT_2___d353 ;

  // register rg_mpie
  always@(MUX_rg_mie_write_1__SEL_1 or
	  write_csr_word or
	  MUX_rg_mie_write_1__SEL_2 or MUX_rg_mcause_write_1__SEL_2 or rg_mie)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_rg_mie_write_1__SEL_1: rg_mpie_D_IN = write_csr_word[7];
      MUX_rg_mie_write_1__SEL_2: rg_mpie_D_IN = 1'd1;
      MUX_rg_mcause_write_1__SEL_2: rg_mpie_D_IN = rg_mie;
      default: rg_mpie_D_IN = 1'b0 /* unspecified value */ ;
    endcase
  end
  assign rg_mpie_EN =
	     EN_write_csr && write_csr_addr == 12'h300 ||
	     EN_upd_on_ret && upd_on_ret_prv == 2'd3 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_mpp
  always@(MUX_rg_mie_write_1__SEL_2 or
	  MUX_rg_mcause_write_1__SEL_2 or
	  mv_curr_priv or MUX_rg_mpp_write_1__SEL_3 or write_csr_word)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_rg_mie_write_1__SEL_2: rg_mpp_D_IN = 2'd0;
      MUX_rg_mcause_write_1__SEL_2: rg_mpp_D_IN = mv_curr_priv;
      MUX_rg_mpp_write_1__SEL_3: rg_mpp_D_IN = write_csr_word[12:11];
      default: rg_mpp_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign rg_mpp_EN =
	     EN_upd_on_ret && upd_on_ret_prv == 2'd3 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ||
	     MUX_rg_mpp_write_1__SEL_3 ;

  // register rg_mprv
  assign rg_mprv_D_IN = write_csr_word[17] ;
  assign rg_mprv_EN = MUX_rg_mie_write_1__SEL_1 ;

  // register rg_mscratch
  assign rg_mscratch_D_IN = write_csr_word ;
  assign rg_mscratch_EN = EN_write_csr && write_csr_addr == 12'h340 ;

  // register rg_msie
  assign rg_msie_D_IN = write_csr_word[3] ;
  assign rg_msie_EN = EN_write_csr && write_csr_addr == 12'h304 ;

  // register rg_msip
  assign rg_msip_D_IN = clint_msip_intrpt ;
  assign rg_msip_EN = EN_clint_msip ;

  // register rg_mtie
  assign rg_mtie_D_IN = write_csr_word[7] ;
  assign rg_mtie_EN = EN_write_csr && write_csr_addr == 12'h304 ;

  // register rg_mtip
  assign rg_mtip_D_IN = clint_mtip_intrpt ;
  assign rg_mtip_EN = EN_clint_mtip ;

  // register rg_mtval
  assign rg_mtval_D_IN =
	     MUX_rg_mtval_write_1__SEL_1 ? write_csr_word : upd_on_trap_tval ;
  assign rg_mtval_EN =
	     EN_write_csr && write_csr_addr == 12'h343 ||
	     EN_upd_on_trap &&
	     NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 ;

  // register rg_mtvec
  assign rg_mtvec_D_IN = { 32'd0, write_csr_word[31:2] } ;
  assign rg_mtvec_EN = EN_write_csr && write_csr_addr == 12'h305 ;

  // register rg_prv
  assign rg_prv_D_IN =
	     EN_upd_on_ret ?
	       MUX_rg_prv_write_1__VAL_1 :
	       MUX_rg_prv_write_1__VAL_2 ;
  assign rg_prv_EN = EN_upd_on_ret || EN_upd_on_trap ;

  // register rg_ucause
  assign rg_ucause_D_IN =
	     MUX_rg_ucause_write_1__SEL_1 ?
	       upd_on_trap_cause[4:0] :
	       write_csr_word[4:0] ;
  assign rg_ucause_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr && write_csr_addr == 12'h042 ;

  // register rg_ueie
  assign rg_ueie_D_IN = write_csr_word[8] ;
  assign rg_ueie_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h304 || write_csr_addr == 12'h004) ;

  // register rg_uepc
  assign rg_uepc_D_IN =
	     MUX_rg_ucause_write_1__SEL_1 ?
	       upd_on_trap_pc[63:1] :
	       write_csr_word[63:1] ;
  assign rg_uepc_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr && write_csr_addr == 12'h041 ;

  // register rg_uie
  always@(MUX_rg_ucause_write_1__SEL_1 or
	  MUX_rg_uie_write_1__SEL_2 or
	  write_csr_word or MUX_rg_uie_write_1__SEL_3 or rg_upie)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_rg_ucause_write_1__SEL_1: rg_uie_D_IN = 1'd0;
      MUX_rg_uie_write_1__SEL_2: rg_uie_D_IN = write_csr_word[0];
      MUX_rg_uie_write_1__SEL_3: rg_uie_D_IN = rg_upie;
      default: rg_uie_D_IN = 1'b0 /* unspecified value */ ;
    endcase
  end
  assign rg_uie_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr &&
	     (write_csr_addr == 12'h300 || write_csr_addr == 12'h0) ||
	     EN_upd_on_ret && upd_on_ret_prv != 2'd3 ;

  // register rg_uinterrupt
  assign rg_uinterrupt_D_IN =
	     MUX_rg_ucause_write_1__SEL_1 ?
	       upd_on_trap_cause[5] :
	       write_csr_word[63] ;
  assign rg_uinterrupt_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr && write_csr_addr == 12'h042 ;

  // register rg_umode
  assign rg_umode_D_IN = write_csr_word[1:0] ;
  assign rg_umode_EN =
	     EN_write_csr && write_csr_addr == 12'h005 &&
	     write_csr_word_BITS_1_TO_0_52_ULT_2___d353 ;

  // register rg_upie
  always@(MUX_rg_ucause_write_1__SEL_1 or
	  rg_uie or
	  MUX_rg_uie_write_1__SEL_2 or
	  write_csr_word or MUX_rg_uie_write_1__SEL_3)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_rg_ucause_write_1__SEL_1: rg_upie_D_IN = rg_uie;
      MUX_rg_uie_write_1__SEL_2: rg_upie_D_IN = write_csr_word[4];
      MUX_rg_uie_write_1__SEL_3: rg_upie_D_IN = 1'd1;
      default: rg_upie_D_IN = 1'b0 /* unspecified value */ ;
    endcase
  end
  assign rg_upie_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr &&
	     (write_csr_addr == 12'h300 || write_csr_addr == 12'h0) ||
	     EN_upd_on_ret && upd_on_ret_prv != 2'd3 ;

  // register rg_uscratch
  assign rg_uscratch_D_IN = write_csr_word ;
  assign rg_uscratch_EN = EN_write_csr && write_csr_addr == 12'h040 ;

  // register rg_usie
  assign rg_usie_D_IN = write_csr_word[0] ;
  assign rg_usie_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h304 || write_csr_addr == 12'h004) ;

  // register rg_usip
  assign rg_usip_D_IN = write_csr_word[0] ;
  assign rg_usip_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h344 || write_csr_addr == 12'h044) &&
	     misa_n ;

  // register rg_utie
  assign rg_utie_D_IN = write_csr_word[4] ;
  assign rg_utie_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h304 || write_csr_addr == 12'h004) ;

  // register rg_utip
  assign rg_utip_D_IN = write_csr_word[4] ;
  assign rg_utip_EN = EN_write_csr && write_csr_addr == 12'h344 && misa_n ;

  // register rg_utval
  assign rg_utval_D_IN =
	     MUX_rg_ucause_write_1__SEL_1 ?
	       upd_on_trap_tval :
	       write_csr_word ;
  assign rg_utval_EN =
	     EN_upd_on_trap &&
	     rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 ||
	     EN_write_csr && write_csr_addr == 12'h043 ;

  // register rg_utvec
  assign rg_utvec_D_IN = { 32'd0, write_csr_word[31:2] } ;
  assign rg_utvec_EN = EN_write_csr && write_csr_addr == 12'h005 ;

  // register soft_ueip
  assign soft_ueip_D_IN = write_csr_word[8] ;
  assign soft_ueip_EN =
	     EN_write_csr &&
	     (write_csr_addr == 12'h344 || write_csr_addr == 12'h044) &&
	     misa_n ;

  // register trigger_index
  assign trigger_index_D_IN = write_csr_word[0] ;
  assign trigger_index_EN = EN_write_csr && write_csr_addr == 12'h7A0 ;

  // register v_pmp_addr_0
  assign v_pmp_addr_0_D_IN = write_csr_word[29:0] ;
  assign v_pmp_addr_0_EN =
	     EN_write_csr && write_csr_addr == 12'h3B0 && !v_pmp_cfg_0[7] ;

  // register v_pmp_addr_1
  assign v_pmp_addr_1_D_IN = write_csr_word[29:0] ;
  assign v_pmp_addr_1_EN =
	     EN_write_csr && write_csr_addr == 12'h3B1 && !v_pmp_cfg_1[7] ;

  // register v_pmp_addr_2
  assign v_pmp_addr_2_D_IN = write_csr_word[29:0] ;
  assign v_pmp_addr_2_EN =
	     EN_write_csr && write_csr_addr == 12'h3B2 && !v_pmp_cfg_2[7] ;

  // register v_pmp_addr_3
  assign v_pmp_addr_3_D_IN = write_csr_word[29:0] ;
  assign v_pmp_addr_3_EN =
	     EN_write_csr && write_csr_addr == 12'h3B3 && !v_pmp_cfg_3[7] ;

  // register v_pmp_cfg_0
  assign v_pmp_cfg_0_D_IN = write_csr_word[7:0] ;
  assign v_pmp_cfg_0_EN =
	     EN_write_csr && write_csr_addr == 12'h3A0 && !v_pmp_cfg_0[7] ;

  // register v_pmp_cfg_1
  assign v_pmp_cfg_1_D_IN = write_csr_word[15:8] ;
  assign v_pmp_cfg_1_EN =
	     EN_write_csr && write_csr_addr == 12'h3A0 && !v_pmp_cfg_1[7] ;

  // register v_pmp_cfg_2
  assign v_pmp_cfg_2_D_IN = write_csr_word[23:16] ;
  assign v_pmp_cfg_2_EN =
	     EN_write_csr && write_csr_addr == 12'h3A0 && !v_pmp_cfg_2[7] ;

  // register v_pmp_cfg_3
  assign v_pmp_cfg_3_D_IN = write_csr_word[31:24] ;
  assign v_pmp_cfg_3_EN =
	     EN_write_csr && write_csr_addr == 12'h3A0 && !v_pmp_cfg_3[7] ;

  // register v_tinfo_0
  assign v_tinfo_0_D_IN = 64'h0 ;
  assign v_tinfo_0_EN = 1'b0 ;

  // register v_tinfo_1
  assign v_tinfo_1_D_IN = 64'h0 ;
  assign v_tinfo_1_EN = 1'b0 ;

  // register v_trig_tdata1_0
  assign v_trig_tdata1_0_D_IN = v_trig_tdata1_1_D_IN ;
  assign v_trig_tdata1_0_EN =
	     EN_write_csr && trigger_index == 1'd0 &&
	     write_csr_addr == 12'h7A1 ;

  // register v_trig_tdata1_1
  always@(write_csr_word or x__h9596 or x__h9759)
  begin
    case (write_csr_word[63:60])
      4'd2:
	  v_trig_tdata1_1_D_IN =
	      { 2'd0,
		write_csr_word[0],
		write_csr_word[1],
		write_csr_word[2],
		write_csr_word[3],
		write_csr_word[6],
		x__h9596,
		write_csr_word[11],
		write_csr_word[15:12],
		x__h9759,
		write_csr_word[19:18] };
      4'd4:
	  v_trig_tdata1_1_D_IN =
	      { 2'd1,
		11'b01010101010 /* unspecified value */ ,
		write_csr_word[5:0],
		write_csr_word[6],
		write_csr_word[9:8] };
      4'd5:
	  v_trig_tdata1_1_D_IN =
	      { 2'd2,
		11'b01010101010 /* unspecified value */ ,
		write_csr_word[5:0],
		write_csr_word[6],
		write_csr_word[9:8] };
      default: v_trig_tdata1_1_D_IN =
		   { 2'd3,
		     20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  assign v_trig_tdata1_1_EN =
	     EN_write_csr && trigger_index == 1'd1 &&
	     write_csr_addr == 12'h7A1 ;

  // register v_trig_tdata2_0
  assign v_trig_tdata2_0_D_IN = write_csr_word ;
  assign v_trig_tdata2_0_EN =
	     EN_write_csr && trigger_index == 1'd0 &&
	     write_csr_addr == 12'h7A2 ;

  // register v_trig_tdata2_1
  assign v_trig_tdata2_1_D_IN = write_csr_word ;
  assign v_trig_tdata2_1_EN =
	     EN_write_csr && trigger_index == 1'd1 &&
	     write_csr_addr == 12'h7A2 ;

  // register v_trig_tdata3_0
  assign v_trig_tdata3_0_D_IN = write_csr_word[50] ;
  assign v_trig_tdata3_0_EN =
	     EN_write_csr && trigger_index == 1'd0 &&
	     write_csr_addr == 12'h7A3 ;

  // register v_trig_tdata3_1
  assign v_trig_tdata3_1_D_IN = write_csr_word[50] ;
  assign v_trig_tdata3_1_EN =
	     EN_write_csr && trigger_index == 1'd1 &&
	     write_csr_addr == 12'h7A3 ;

  // remaining internal signals
  assign IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d117 =
	     CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q20 ?
	       { 4'd5,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45,
		 49'd0,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d109 } :
	       64'd0 ;
  assign IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d118 =
	     CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q21 ?
	       { 4'd4,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45,
		 49'd0,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d109 } :
	       IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d117 ;
  assign IF_rg_mode_77_EQ_1_10_AND_upd_on_trap_cause_BI_ETC___d713 =
	     (rg_mode == 2'd1 && upd_on_trap_cause[5]) ?
	       rg_mtvec + { 57'd0, upd_on_trap_cause[4:0] } :
	       rg_mtvec ;
  assign IF_rg_umode_75_EQ_1_05_AND_upd_on_trap_cause_B_ETC___d709 =
	     (rg_umode == 2'd1 && upd_on_trap_cause[5]) ?
	       rg_utvec + { 57'd0, upd_on_trap_cause[4:0] } :
	       rg_utvec ;
  assign IF_upd_on_ret_prv_EQ_3_41_THEN_IF_misa_c_83_TH_ETC___d652 =
	     (upd_on_ret_prv == 2'd3) ?
	       (misa_c ? rg_mepc : result__h10415) :
	       (misa_c ? rg_uepc : result__h10268) ;
  assign NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691 =
	     !rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d669 &&
	     !rg_medeleg_u1_56_CONCAT_0_CONCAT_rg_medeleg_m2_ETC___d673 ||
	     rg_prv == 2'd3 ||
	     !misa_n ;
  assign SEL_ARR_v_trig_tdata1_0_4_BITS_14_TO_11_4_v_tr_ETC___d90 =
	     { CASE_trigger_index_0_v_trig_tdata1_0_BITS_14_T_ETC__q15,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_15_1__ETC__q16,
	       2'd0,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_16_1__ETC__q17,
	       SEL_ARR_v_trig_tdata1_0_4_BIT_17_6_v_trig_tdat_ETC___d88 } ;
  assign SEL_ARR_v_trig_tdata1_0_4_BITS_9_TO_6_6_v_trig_ETC___d91 =
	     { CASE_trigger_index_0_v_trig_tdata1_0_BITS_9_TO_ETC__q18,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_10_1__ETC__q19,
	       SEL_ARR_v_trig_tdata1_0_4_BITS_14_TO_11_4_v_tr_ETC___d90 } ;
  assign SEL_ARR_v_trig_tdata1_0_4_BIT_17_6_v_trig_tdat_ETC___d88 =
	     { CASE_trigger_index_0_v_trig_tdata1_0_BIT_17_1__ETC__q12,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_18_1__ETC__q13,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_19_1__ETC__q14 } ;
  assign SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d109 =
	     { SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d54,
	       2'd0,
	       CASE_trigger_index_0_v_trig_tdata1_0_BIT_2_1_v_ETC__q10,
	       CASE_trigger_index_0_v_trig_tdata1_0_BITS_8_TO_ETC__q11 } ;
  assign _0_CONCAT_rg_utie_82_AND_misa_n_45_AND_rg_utip__ETC___d738 =
	     { 2'd0,
	       rg_utie & misa_n_45_AND_rg_utip_49___d239,
	       rg_msie & rg_msip,
	       2'd0,
	       rg_usie & misa_n_45_AND_rg_usip_54___d240 } ;
  assign _theResult_____2__h3288 = read_csr ;
  assign data___1__h3506 =
	     { 13'd0,
	       CASE_trigger_index_0_v_trig_tdata3_0_1_v_trig__ETC__q7,
	       50'd0 } ;
  assign data___1__h3703 =
	     CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q22 ?
	       { 4'd2,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45,
		 36'd0,
		 SEL_ARR_v_trig_tdata1_0_4_BITS_5_TO_2_6_v_trig_ETC___d49[3:2],
		 1'b0,
		 SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d54,
		 1'b0,
		 SEL_ARR_v_trig_tdata1_0_4_BITS_5_TO_2_6_v_trig_ETC___d49[1:0],
		 SEL_ARR_v_trig_tdata1_0_4_BITS_9_TO_6_6_v_trig_ETC___d91 } :
	       IF_SEL_ARR_v_trig_tdata1_0_4_BITS_21_TO_20_5_E_ETC___d118 ;
  assign data___1__h4095 = { 63'd0, trigger_index } ;
  assign data___1__h4119 = { 56'd0, x__h4122 } ;
  assign data___1__h4126 = { 61'd0, frm } ;
  assign data___1__h4131 = { 59'd0, fflags } ;
  assign data___1__h4147 =
	     { 52'd0,
	       rg_meip,
	       2'd0,
	       x__h4161 & misa_n,
	       rg_mtip,
	       2'd0,
	       x__h4195 & misa_n,
	       rg_msip,
	       2'd0,
	       x__h4223 & misa_n } ;
  assign data___1__h4262 = { rg_uinterrupt, 58'd0, rg_ucause } ;
  assign data___1__h4273 = { rg_uepc, 1'b0 } ;
  assign data___1__h4282 = { rg_utvec, rg_umode } ;
  assign data___1__h4287 =
	     { 52'd0,
	       rg_meie,
	       2'd0,
	       rg_mideleg[8] & rg_ueie,
	       rg_mtie,
	       2'd0,
	       rg_mideleg[4] & rg_utie,
	       rg_msie,
	       2'd0,
	       rg_mideleg[0] & rg_usie } ;
  assign data___1__h4391 =
	     { r__h4396, 48'd262144, fs, 8'd0, rg_upie, 3'd0, rg_uie } ;
  assign data___1__h4458 = { 34'd0, v_pmp_addr_3 } ;
  assign data___1__h4603 = { 34'd0, v_pmp_addr_2 } ;
  assign data___1__h4620 = { 34'd0, v_pmp_addr_1 } ;
  assign data___1__h4637 = { 34'd0, v_pmp_addr_0 } ;
  assign data___1__h4730 =
	     { 32'd0, v_pmp_cfg_3, v_pmp_cfg_2, v_pmp_cfg_1, v_pmp_cfg_0 } ;
  assign data___1__h5125 = { 61'd0, rg_mcounteren } ;
  assign data___1__h5131 = { rg_minterrupt, 58'd0, rg_mcause } ;
  assign data___1__h5145 = { rg_mepc, 1'b0 } ;
  assign data___1__h5155 =
	     { 52'd0,
	       rg_meip,
	       2'd0,
	       misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238,
	       rg_mtip,
	       2'd0,
	       misa_n_45_AND_rg_utip_49___d239,
	       rg_msip,
	       2'd0,
	       misa_n_45_AND_rg_usip_54___d240 } ;
  assign data___1__h5188 =
	     { 52'd0,
	       rg_meie,
	       2'd0,
	       misa_n_45_AND_rg_ueie_79___d247,
	       rg_mtie,
	       2'd0,
	       misa_n_45_AND_rg_utie_82___d248,
	       rg_msie,
	       2'd0,
	       misa_n_45_AND_rg_usie_85___d249 } ;
  assign data___1__h5221 =
	     { 48'd0,
	       rg_medeleg_u1,
	       1'd0,
	       rg_medeleg_m2,
	       2'd0,
	       rg_medeleg_l10 } ;
  assign data___1__h5230 = { 52'd0, rg_mideleg } ;
  assign data___1__h5232 =
	     { r__h4396,
	       45'd163840,
	       rg_mprv,
	       2'd0,
	       fs,
	       rg_mpp,
	       3'd0,
	       rg_mpie,
	       2'd0,
	       rg_upie,
	       rg_mie,
	       2'd0,
	       rg_uie } ;
  assign data___1__h5260 = { rg_mtvec, rg_mode } ;
  assign misa__h262 =
	     { 5'd0,
	       misa_u,
	       6'd16,
	       misa_n,
	       misa_m,
	       3'd0,
	       misa_i,
	       5'd0,
	       misa_c,
	       1'd0,
	       misa_a } ;
  assign misa_n_45_AND_rg_ueie_79___d247 = misa_n & rg_ueie ;
  assign misa_n_45_AND_rg_usie_85___d249 = misa_n & rg_usie ;
  assign misa_n_45_AND_rg_usip_54___d240 = misa_n & rg_usip ;
  assign misa_n_45_AND_rg_utie_82___d248 = misa_n & rg_utie ;
  assign misa_n_45_AND_rg_utip_49___d239 = misa_n & rg_utip ;
  assign misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238 =
	     misa_n & y__h4164 ;
  assign mv_csr_decode_csr_mstatus__h15074 = csr_mstatus ;
  assign r__h4396 = fs == 2'b11 ;
  assign result__h10268 = { rg_uepc[62:1], 1'd0 } ;
  assign result__h10415 = { rg_mepc[62:1], 1'd0 } ;
  assign rg_medeleg_u1_56_CONCAT_0_CONCAT_rg_medeleg_m2_ETC___d673 =
	     rg_medeleg_u1_CONCAT_0_CONCAT_rg_medeleg_m2_CO_ETC__q9[0] &
	     ~upd_on_trap_cause[5] ;
  assign rg_medeleg_u1_CONCAT_0_CONCAT_rg_medeleg_m2_CO_ETC__q9 =
	     { rg_medeleg_u1, 1'd0, rg_medeleg_m2, 2'd0, rg_medeleg_l10 } >>
	     upd_on_trap_cause[4:0] ;
  assign rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d669 =
	     rg_mideleg_SRL_upd_on_trap_cause_BITS_4_TO_0__q8[0] &
	     upd_on_trap_cause[5] ;
  assign rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694 =
	     (rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d669 ||
	      rg_medeleg_u1_56_CONCAT_0_CONCAT_rg_medeleg_m2_ETC___d673) &&
	     rg_prv != 2'd3 &&
	     misa_n ;
  assign rg_mideleg_SRL_upd_on_trap_cause_BITS_4_TO_0__q8 =
	     rg_mideleg >> upd_on_trap_cause[4:0] ;
  assign rg_ueie_79_AND_misa_n_45_AND_soft_ueip_41_OR_e_ETC___d739 =
	     { rg_ueie & misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238,
	       rg_mtie & rg_mtip,
	       _0_CONCAT_rg_utie_82_AND_misa_n_45_AND_rg_utip__ETC___d738 } ;
  assign write_csr_addr_EQ_0x1_35_AND_NOT_fflags_25_EQ__ETC___d453 =
	     write_csr_addr == 12'h001 && fflags != write_csr_word[4:0] ||
	     write_csr_addr != 12'h001 &&
	     write_csr_addr_EQ_0x2_41_AND_NOT_frm_24_EQ_wri_ETC___d451 ;
  assign write_csr_addr_EQ_0x2_41_AND_NOT_frm_24_EQ_wri_ETC___d451 =
	     write_csr_addr == 12'h002 && frm != write_csr_word[2:0] ||
	     write_csr_addr == 12'h003 && x__h4122 != write_csr_word[7:0] ;
  assign write_csr_word_BITS_1_TO_0_52_ULT_2___d353 =
	     write_csr_word[1:0] < 2'd2 ;
  assign x__h14812 = mv_curr_priv ;
  assign x__h15117 =
	     { rg_meie,
	       2'd0,
	       rg_ueie,
	       rg_mtie,
	       2'd0,
	       rg_utie,
	       rg_msie,
	       2'd0,
	       rg_usie } ;
  assign x__h15129 =
	     { 3'd0,
	       misa_n_45_AND_soft_ueip_41_OR_ext_ueip_42_43___d238,
	       3'd0,
	       misa_n_45_AND_rg_utip_49___d239,
	       3'd0,
	       misa_n_45_AND_rg_usip_54___d240 } ;
  assign x__h15156 =
	     { 3'd0,
	       misa_n_45_AND_rg_ueie_79___d247,
	       3'd0,
	       misa_n_45_AND_rg_utie_82___d248,
	       3'd0,
	       misa_n_45_AND_rg_usie_85___d249 } ;
  assign x__h15339 =
	     { rg_meie & rg_meip,
	       2'd0,
	       rg_ueie_79_AND_misa_n_45_AND_soft_ueip_41_OR_e_ETC___d739 } ;
  assign x__h4122 = { frm, fflags } ;
  assign x__h4161 = rg_mideleg[8] & y__h4164 ;
  assign x__h4195 = rg_mideleg[4] & rg_utip ;
  assign x__h4223 = rg_mideleg[0] & rg_usip ;
  assign x__h9596 =
	     (!write_csr_word[19] &&
	      (write_csr_word[10:7] == 4'd0 || write_csr_word[10:7] == 4'd2 ||
	       write_csr_word[10:7] == 4'd3)) ?
	       write_csr_word[10:7] :
	       4'd0 ;
  assign x__h9759 = { write_csr_word[22:21], write_csr_word[17:16] } ;
  assign y__h4164 = soft_ueip | ext_ueip ;
  always@(v_trig_tdata1_1)
  begin
    case (v_trig_tdata1_1[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_v_trig_tdata1_1_BITS_21_TO_20_0_v_trig_td_ETC__q1 =
	      v_trig_tdata1_1;
      2'd3:
	  CASE_v_trig_tdata1_1_BITS_21_TO_20_0_v_trig_td_ETC__q1 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(v_trig_tdata1_0)
  begin
    case (v_trig_tdata1_0[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_v_trig_tdata1_0_BITS_21_TO_20_0_v_trig_td_ETC__q2 =
	      v_trig_tdata1_0;
      2'd3:
	  CASE_v_trig_tdata1_0_BITS_21_TO_20_0_v_trig_td_ETC__q2 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(v_trig_tdata1_1)
  begin
    case (v_trig_tdata1_1[21:20])
      2'd1, 2'd2:
	  CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q3 =
	      v_trig_tdata1_1[1];
      default: CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q3 =
		   v_trig_tdata1_1[21:20] == 2'd0 && v_trig_tdata1_1[15];
    endcase
  end
  always@(v_trig_tdata1_1)
  begin
    case (v_trig_tdata1_1[21:20])
      2'd1, 2'd2:
	  CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q4 =
	      v_trig_tdata1_1[2];
      default: CASE_v_trig_tdata1_1_BITS_21_TO_20_1_v_trig_td_ETC__q4 =
		   v_trig_tdata1_1[21:20] == 2'd0 && v_trig_tdata1_1[16];
    endcase
  end
  always@(v_trig_tdata1_0)
  begin
    case (v_trig_tdata1_0[21:20])
      2'd1, 2'd2:
	  CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q5 =
	      v_trig_tdata1_0[1];
      default: CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q5 =
		   v_trig_tdata1_0[21:20] == 2'd0 && v_trig_tdata1_0[15];
    endcase
  end
  always@(v_trig_tdata1_0)
  begin
    case (v_trig_tdata1_0[21:20])
      2'd1, 2'd2:
	  CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q6 =
	      v_trig_tdata1_0[2];
      default: CASE_v_trig_tdata1_0_BITS_21_TO_20_1_v_trig_td_ETC__q6 =
		   v_trig_tdata1_0[21:20] == 2'd0 && v_trig_tdata1_0[16];
    endcase
  end
  always@(trigger_index or v_tinfo_0 or v_tinfo_1)
  begin
    case (trigger_index)
      1'd0: data___1__h3415 = v_tinfo_0;
      1'd1: data___1__h3415 = v_tinfo_1;
    endcase
  end
  always@(trigger_index or v_trig_tdata3_0 or v_trig_tdata3_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata3_0_1_v_trig__ETC__q7 =
	      v_trig_tdata3_0;
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata3_0_1_v_trig__ETC__q7 =
	      v_trig_tdata3_1;
    endcase
  end
  always@(trigger_index or v_trig_tdata2_0 or v_trig_tdata2_1)
  begin
    case (trigger_index)
      1'd0: data___1__h3613 = v_trig_tdata2_0;
      1'd1: data___1__h3613 = v_trig_tdata2_1;
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  SEL_ARR_v_trig_tdata1_0_4_BITS_5_TO_2_6_v_trig_ETC___d49 =
	      v_trig_tdata1_0[5:2];
      1'd1:
	  SEL_ARR_v_trig_tdata1_0_4_BITS_5_TO_2_6_v_trig_ETC___d49 =
	      v_trig_tdata1_1[5:2];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45 =
	      v_trig_tdata1_0[0];
      1'd1:
	  SEL_ARR_v_trig_tdata1_0_4_BIT_0_2_v_trig_tdata_ETC___d45 =
	      v_trig_tdata1_1[0];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d54 =
	      v_trig_tdata1_0[1];
      1'd1:
	  SEL_ARR_v_trig_tdata1_0_4_BIT_1_1_v_trig_tdata_ETC___d54 =
	      v_trig_tdata1_1[1];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_2_1_v_ETC__q10 =
	      v_trig_tdata1_0[2];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_2_1_v_ETC__q10 =
	      v_trig_tdata1_1[2];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_8_TO_ETC__q11 =
	      v_trig_tdata1_0[8:3];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_8_TO_ETC__q11 =
	      v_trig_tdata1_1[8:3];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_17_1__ETC__q12 =
	      v_trig_tdata1_0[17];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_17_1__ETC__q12 =
	      v_trig_tdata1_1[17];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_18_1__ETC__q13 =
	      v_trig_tdata1_0[18];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_18_1__ETC__q13 =
	      v_trig_tdata1_1[18];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_19_1__ETC__q14 =
	      v_trig_tdata1_0[19];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_19_1__ETC__q14 =
	      v_trig_tdata1_1[19];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_14_T_ETC__q15 =
	      v_trig_tdata1_0[14:11];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_14_T_ETC__q15 =
	      v_trig_tdata1_1[14:11];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_15_1__ETC__q16 =
	      v_trig_tdata1_0[15];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_15_1__ETC__q16 =
	      v_trig_tdata1_1[15];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_16_1__ETC__q17 =
	      v_trig_tdata1_0[16];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_16_1__ETC__q17 =
	      v_trig_tdata1_1[16];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_9_TO_ETC__q18 =
	      v_trig_tdata1_0[9:6];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_9_TO_ETC__q18 =
	      v_trig_tdata1_1[9:6];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_10_1__ETC__q19 =
	      v_trig_tdata1_0[10];
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BIT_10_1__ETC__q19 =
	      v_trig_tdata1_1[10];
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q20 =
	      v_trig_tdata1_0[21:20] == 2'd2;
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q20 =
	      v_trig_tdata1_1[21:20] == 2'd2;
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q21 =
	      v_trig_tdata1_0[21:20] == 2'd1;
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q21 =
	      v_trig_tdata1_1[21:20] == 2'd1;
    endcase
  end
  always@(trigger_index or v_trig_tdata1_0 or v_trig_tdata1_1)
  begin
    case (trigger_index)
      1'd0:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q22 =
	      v_trig_tdata1_0[21:20] == 2'd0;
      1'd1:
	  CASE_trigger_index_0_v_trig_tdata1_0_BITS_21_T_ETC__q22 =
	      v_trig_tdata1_1[21:20] == 2'd0;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        ext_ueip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	fflags <= `BSV_ASSIGNMENT_DELAY 5'd0;
	frm <= `BSV_ASSIGNMENT_DELAY 3'd0;
	fs <= `BSV_ASSIGNMENT_DELAY 2'd0;
	mcycle <= `BSV_ASSIGNMENT_DELAY 64'd0;
	minstret <= `BSV_ASSIGNMENT_DELAY 64'd0;
	misa_a <= `BSV_ASSIGNMENT_DELAY 1'd1;
	misa_c <= `BSV_ASSIGNMENT_DELAY 1'd1;
	misa_i <= `BSV_ASSIGNMENT_DELAY 1'd1;
	misa_m <= `BSV_ASSIGNMENT_DELAY 1'd1;
	misa_n <= `BSV_ASSIGNMENT_DELAY 1'd0;
	misa_u <= `BSV_ASSIGNMENT_DELAY 1'd1;
	rg_clint_mtime <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_mcause <= `BSV_ASSIGNMENT_DELAY 5'd0;
	rg_mcounteren <= `BSV_ASSIGNMENT_DELAY 3'd0;
	rg_medeleg_l10 <= `BSV_ASSIGNMENT_DELAY 10'd0;
	rg_medeleg_m2 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	rg_medeleg_u1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_meie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_meip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mepc <= `BSV_ASSIGNMENT_DELAY 63'd0;
	rg_mideleg <= `BSV_ASSIGNMENT_DELAY 12'd0;
	rg_mie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_minterrupt <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mode <= `BSV_ASSIGNMENT_DELAY 2'd0;
	rg_mpie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mpp <= `BSV_ASSIGNMENT_DELAY 2'b0;
	rg_mprv <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mscratch <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_msie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_msip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mtie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mtip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_mtval <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_mtvec <= `BSV_ASSIGNMENT_DELAY 62'd0;
	rg_prv <= `BSV_ASSIGNMENT_DELAY 2'd3;
	rg_ucause <= `BSV_ASSIGNMENT_DELAY 5'd0;
	rg_ueie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_uepc <= `BSV_ASSIGNMENT_DELAY 63'd0;
	rg_uie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_uinterrupt <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_umode <= `BSV_ASSIGNMENT_DELAY 2'd0;
	rg_upie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_uscratch <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_usie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_usip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_utie <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_utip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_utval <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_utvec <= `BSV_ASSIGNMENT_DELAY 62'd0;
	soft_ueip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	trigger_index <= `BSV_ASSIGNMENT_DELAY 1'd0;
	v_pmp_addr_0 <= `BSV_ASSIGNMENT_DELAY 30'd0;
	v_pmp_addr_1 <= `BSV_ASSIGNMENT_DELAY 30'd0;
	v_pmp_addr_2 <= `BSV_ASSIGNMENT_DELAY 30'd0;
	v_pmp_addr_3 <= `BSV_ASSIGNMENT_DELAY 30'd0;
	v_pmp_cfg_0 <= `BSV_ASSIGNMENT_DELAY 8'd0;
	v_pmp_cfg_1 <= `BSV_ASSIGNMENT_DELAY 8'd0;
	v_pmp_cfg_2 <= `BSV_ASSIGNMENT_DELAY 8'd0;
	v_pmp_cfg_3 <= `BSV_ASSIGNMENT_DELAY 8'd0;
	v_tinfo_0 <= `BSV_ASSIGNMENT_DELAY 64'd52;
	v_tinfo_1 <= `BSV_ASSIGNMENT_DELAY 64'd52;
	v_trig_tdata1_0 <= `BSV_ASSIGNMENT_DELAY
	    { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
	v_trig_tdata1_1 <= `BSV_ASSIGNMENT_DELAY
	    { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
	v_trig_tdata2_0 <= `BSV_ASSIGNMENT_DELAY 64'd0;
	v_trig_tdata2_1 <= `BSV_ASSIGNMENT_DELAY 64'd0;
	v_trig_tdata3_0 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	v_trig_tdata3_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (ext_ueip_EN) ext_ueip <= `BSV_ASSIGNMENT_DELAY ext_ueip_D_IN;
	if (fflags_EN) fflags <= `BSV_ASSIGNMENT_DELAY fflags_D_IN;
	if (frm_EN) frm <= `BSV_ASSIGNMENT_DELAY frm_D_IN;
	if (fs_EN) fs <= `BSV_ASSIGNMENT_DELAY fs_D_IN;
	if (mcycle_EN) mcycle <= `BSV_ASSIGNMENT_DELAY mcycle_D_IN;
	if (minstret_EN) minstret <= `BSV_ASSIGNMENT_DELAY minstret_D_IN;
	if (misa_a_EN) misa_a <= `BSV_ASSIGNMENT_DELAY misa_a_D_IN;
	if (misa_c_EN) misa_c <= `BSV_ASSIGNMENT_DELAY misa_c_D_IN;
	if (misa_i_EN) misa_i <= `BSV_ASSIGNMENT_DELAY misa_i_D_IN;
	if (misa_m_EN) misa_m <= `BSV_ASSIGNMENT_DELAY misa_m_D_IN;
	if (misa_n_EN) misa_n <= `BSV_ASSIGNMENT_DELAY misa_n_D_IN;
	if (misa_u_EN) misa_u <= `BSV_ASSIGNMENT_DELAY misa_u_D_IN;
	if (rg_clint_mtime_EN)
	  rg_clint_mtime <= `BSV_ASSIGNMENT_DELAY rg_clint_mtime_D_IN;
	if (rg_mcause_EN) rg_mcause <= `BSV_ASSIGNMENT_DELAY rg_mcause_D_IN;
	if (rg_mcounteren_EN)
	  rg_mcounteren <= `BSV_ASSIGNMENT_DELAY rg_mcounteren_D_IN;
	if (rg_medeleg_l10_EN)
	  rg_medeleg_l10 <= `BSV_ASSIGNMENT_DELAY rg_medeleg_l10_D_IN;
	if (rg_medeleg_m2_EN)
	  rg_medeleg_m2 <= `BSV_ASSIGNMENT_DELAY rg_medeleg_m2_D_IN;
	if (rg_medeleg_u1_EN)
	  rg_medeleg_u1 <= `BSV_ASSIGNMENT_DELAY rg_medeleg_u1_D_IN;
	if (rg_meie_EN) rg_meie <= `BSV_ASSIGNMENT_DELAY rg_meie_D_IN;
	if (rg_meip_EN) rg_meip <= `BSV_ASSIGNMENT_DELAY rg_meip_D_IN;
	if (rg_mepc_EN) rg_mepc <= `BSV_ASSIGNMENT_DELAY rg_mepc_D_IN;
	if (rg_mideleg_EN)
	  rg_mideleg <= `BSV_ASSIGNMENT_DELAY rg_mideleg_D_IN;
	if (rg_mie_EN) rg_mie <= `BSV_ASSIGNMENT_DELAY rg_mie_D_IN;
	if (rg_minterrupt_EN)
	  rg_minterrupt <= `BSV_ASSIGNMENT_DELAY rg_minterrupt_D_IN;
	if (rg_mode_EN) rg_mode <= `BSV_ASSIGNMENT_DELAY rg_mode_D_IN;
	if (rg_mpie_EN) rg_mpie <= `BSV_ASSIGNMENT_DELAY rg_mpie_D_IN;
	if (rg_mpp_EN) rg_mpp <= `BSV_ASSIGNMENT_DELAY rg_mpp_D_IN;
	if (rg_mprv_EN) rg_mprv <= `BSV_ASSIGNMENT_DELAY rg_mprv_D_IN;
	if (rg_mscratch_EN)
	  rg_mscratch <= `BSV_ASSIGNMENT_DELAY rg_mscratch_D_IN;
	if (rg_msie_EN) rg_msie <= `BSV_ASSIGNMENT_DELAY rg_msie_D_IN;
	if (rg_msip_EN) rg_msip <= `BSV_ASSIGNMENT_DELAY rg_msip_D_IN;
	if (rg_mtie_EN) rg_mtie <= `BSV_ASSIGNMENT_DELAY rg_mtie_D_IN;
	if (rg_mtip_EN) rg_mtip <= `BSV_ASSIGNMENT_DELAY rg_mtip_D_IN;
	if (rg_mtval_EN) rg_mtval <= `BSV_ASSIGNMENT_DELAY rg_mtval_D_IN;
	if (rg_mtvec_EN) rg_mtvec <= `BSV_ASSIGNMENT_DELAY rg_mtvec_D_IN;
	if (rg_prv_EN) rg_prv <= `BSV_ASSIGNMENT_DELAY rg_prv_D_IN;
	if (rg_ucause_EN) rg_ucause <= `BSV_ASSIGNMENT_DELAY rg_ucause_D_IN;
	if (rg_ueie_EN) rg_ueie <= `BSV_ASSIGNMENT_DELAY rg_ueie_D_IN;
	if (rg_uepc_EN) rg_uepc <= `BSV_ASSIGNMENT_DELAY rg_uepc_D_IN;
	if (rg_uie_EN) rg_uie <= `BSV_ASSIGNMENT_DELAY rg_uie_D_IN;
	if (rg_uinterrupt_EN)
	  rg_uinterrupt <= `BSV_ASSIGNMENT_DELAY rg_uinterrupt_D_IN;
	if (rg_umode_EN) rg_umode <= `BSV_ASSIGNMENT_DELAY rg_umode_D_IN;
	if (rg_upie_EN) rg_upie <= `BSV_ASSIGNMENT_DELAY rg_upie_D_IN;
	if (rg_uscratch_EN)
	  rg_uscratch <= `BSV_ASSIGNMENT_DELAY rg_uscratch_D_IN;
	if (rg_usie_EN) rg_usie <= `BSV_ASSIGNMENT_DELAY rg_usie_D_IN;
	if (rg_usip_EN) rg_usip <= `BSV_ASSIGNMENT_DELAY rg_usip_D_IN;
	if (rg_utie_EN) rg_utie <= `BSV_ASSIGNMENT_DELAY rg_utie_D_IN;
	if (rg_utip_EN) rg_utip <= `BSV_ASSIGNMENT_DELAY rg_utip_D_IN;
	if (rg_utval_EN) rg_utval <= `BSV_ASSIGNMENT_DELAY rg_utval_D_IN;
	if (rg_utvec_EN) rg_utvec <= `BSV_ASSIGNMENT_DELAY rg_utvec_D_IN;
	if (soft_ueip_EN) soft_ueip <= `BSV_ASSIGNMENT_DELAY soft_ueip_D_IN;
	if (trigger_index_EN)
	  trigger_index <= `BSV_ASSIGNMENT_DELAY trigger_index_D_IN;
	if (v_pmp_addr_0_EN)
	  v_pmp_addr_0 <= `BSV_ASSIGNMENT_DELAY v_pmp_addr_0_D_IN;
	if (v_pmp_addr_1_EN)
	  v_pmp_addr_1 <= `BSV_ASSIGNMENT_DELAY v_pmp_addr_1_D_IN;
	if (v_pmp_addr_2_EN)
	  v_pmp_addr_2 <= `BSV_ASSIGNMENT_DELAY v_pmp_addr_2_D_IN;
	if (v_pmp_addr_3_EN)
	  v_pmp_addr_3 <= `BSV_ASSIGNMENT_DELAY v_pmp_addr_3_D_IN;
	if (v_pmp_cfg_0_EN)
	  v_pmp_cfg_0 <= `BSV_ASSIGNMENT_DELAY v_pmp_cfg_0_D_IN;
	if (v_pmp_cfg_1_EN)
	  v_pmp_cfg_1 <= `BSV_ASSIGNMENT_DELAY v_pmp_cfg_1_D_IN;
	if (v_pmp_cfg_2_EN)
	  v_pmp_cfg_2 <= `BSV_ASSIGNMENT_DELAY v_pmp_cfg_2_D_IN;
	if (v_pmp_cfg_3_EN)
	  v_pmp_cfg_3 <= `BSV_ASSIGNMENT_DELAY v_pmp_cfg_3_D_IN;
	if (v_tinfo_0_EN) v_tinfo_0 <= `BSV_ASSIGNMENT_DELAY v_tinfo_0_D_IN;
	if (v_tinfo_1_EN) v_tinfo_1 <= `BSV_ASSIGNMENT_DELAY v_tinfo_1_D_IN;
	if (v_trig_tdata1_0_EN)
	  v_trig_tdata1_0 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata1_0_D_IN;
	if (v_trig_tdata1_1_EN)
	  v_trig_tdata1_1 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata1_1_D_IN;
	if (v_trig_tdata2_0_EN)
	  v_trig_tdata2_0 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata2_0_D_IN;
	if (v_trig_tdata2_1_EN)
	  v_trig_tdata2_1 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata2_1_D_IN;
	if (v_trig_tdata3_0_EN)
	  v_trig_tdata3_0 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata3_0_D_IN;
	if (v_trig_tdata3_1_EN)
	  v_trig_tdata3_1 <= `BSV_ASSIGNMENT_DELAY v_trig_tdata3_1_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    ext_ueip = 1'h0;
    fflags = 5'h0A;
    frm = 3'h2;
    fs = 2'h2;
    mcycle = 64'hAAAAAAAAAAAAAAAA;
    minstret = 64'hAAAAAAAAAAAAAAAA;
    misa_a = 1'h0;
    misa_c = 1'h0;
    misa_i = 1'h0;
    misa_m = 1'h0;
    misa_n = 1'h0;
    misa_u = 1'h0;
    rg_clint_mtime = 64'hAAAAAAAAAAAAAAAA;
    rg_mcause = 5'h0A;
    rg_mcounteren = 3'h2;
    rg_medeleg_l10 = 10'h2AA;
    rg_medeleg_m2 = 2'h2;
    rg_medeleg_u1 = 1'h0;
    rg_meie = 1'h0;
    rg_meip = 1'h0;
    rg_mepc = 63'h2AAAAAAAAAAAAAAA;
    rg_mideleg = 12'hAAA;
    rg_mie = 1'h0;
    rg_minterrupt = 1'h0;
    rg_mode = 2'h2;
    rg_mpie = 1'h0;
    rg_mpp = 2'h2;
    rg_mprv = 1'h0;
    rg_mscratch = 64'hAAAAAAAAAAAAAAAA;
    rg_msie = 1'h0;
    rg_msip = 1'h0;
    rg_mtie = 1'h0;
    rg_mtip = 1'h0;
    rg_mtval = 64'hAAAAAAAAAAAAAAAA;
    rg_mtvec = 62'h2AAAAAAAAAAAAAAA;
    rg_prv = 2'h2;
    rg_ucause = 5'h0A;
    rg_ueie = 1'h0;
    rg_uepc = 63'h2AAAAAAAAAAAAAAA;
    rg_uie = 1'h0;
    rg_uinterrupt = 1'h0;
    rg_umode = 2'h2;
    rg_upie = 1'h0;
    rg_uscratch = 64'hAAAAAAAAAAAAAAAA;
    rg_usie = 1'h0;
    rg_usip = 1'h0;
    rg_utie = 1'h0;
    rg_utip = 1'h0;
    rg_utval = 64'hAAAAAAAAAAAAAAAA;
    rg_utvec = 62'h2AAAAAAAAAAAAAAA;
    soft_ueip = 1'h0;
    trigger_index = 1'h0;
    v_pmp_addr_0 = 30'h2AAAAAAA;
    v_pmp_addr_1 = 30'h2AAAAAAA;
    v_pmp_addr_2 = 30'h2AAAAAAA;
    v_pmp_addr_3 = 30'h2AAAAAAA;
    v_pmp_cfg_0 = 8'hAA;
    v_pmp_cfg_1 = 8'hAA;
    v_pmp_cfg_2 = 8'hAA;
    v_pmp_cfg_3 = 8'hAA;
    v_tinfo_0 = 64'hAAAAAAAAAAAAAAAA;
    v_tinfo_1 = 64'hAAAAAAAAAAAAAAAA;
    v_trig_tdata1_0 = 22'h2AAAAA;
    v_trig_tdata1_1 = 22'h2AAAAA;
    v_trig_tdata2_0 = 64'hAAAAAAAAAAAAAAAA;
    v_trig_tdata2_1 = 64'hAAAAAAAAAAAAAAAA;
    v_trig_tdata3_0 = 1'h0;
    v_trig_tdata3_1 = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d3 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d4 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d5 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  v__h3202 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d3 ||
	   TASK_testplusargs___d4 && TASK_testplusargs___d5))
	$write("[%10d", v__h3202, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d3 ||
	   TASK_testplusargs___d4 && TASK_testplusargs___d5))
	$write("CSRFILE : Read Operation : Addr:%h", read_csr_addr);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d3 ||
	   TASK_testplusargs___d4 && TASK_testplusargs___d5))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d9 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d10 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  TASK_testplusargs___d11 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr)
	begin
	  v__h3355 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d9 ||
	   TASK_testplusargs___d10 && TASK_testplusargs___d11))
	$write("[%10d", v__h3355, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d9 ||
	   TASK_testplusargs___d10 && TASK_testplusargs___d11))
	$write("CSRFILE : Read Operation : Addr:%h Data:%h",
	       read_csr_addr,
	       _theResult_____2__h3288);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_read_csr &&
	  (TASK_testplusargs___d9 ||
	   TASK_testplusargs___d10 && TASK_testplusargs___d11))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr)
	begin
	  TASK_testplusargs___d333 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr)
	begin
	  TASK_testplusargs___d334 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr)
	begin
	  TASK_testplusargs___d335 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr)
	begin
	  v__h5566 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr &&
	  (TASK_testplusargs___d333 ||
	   TASK_testplusargs___d334 && TASK_testplusargs___d335))
	$write("[%10d", v__h5566, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr &&
	  (TASK_testplusargs___d333 ||
	   TASK_testplusargs___d334 && TASK_testplusargs___d335))
	$write("CSRFILE : Write Operation : Addr:%h, word:%h",
	       write_csr_addr,
	       write_csr_word);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_write_csr &&
	  (TASK_testplusargs___d333 ||
	   TASK_testplusargs___d334 && TASK_testplusargs___d335))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d653 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d654 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d655 = $test$plusargs("l2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  v__h10538 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d653 ||
	   TASK_testplusargs___d654 && TASK_testplusargs___d655))
	$write("[%10d", v__h10538, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d653 ||
	   TASK_testplusargs___d654 && TASK_testplusargs___d655))
	$write("CSRFILE : PC:%h Cause:%d misa_s:%b",
	       upd_on_trap_pc,
	       upd_on_trap_cause,
	       1'd1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d653 ||
	   TASK_testplusargs___d654 && TASK_testplusargs___d655))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d659 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d660 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d661 = $test$plusargs("l2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  v__h10688 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d659 ||
	   TASK_testplusargs___d660 && TASK_testplusargs___d661))
	$write("[%10d", v__h10688, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d659 ||
	   TASK_testplusargs___d660 && TASK_testplusargs___d661))
	$write("CSRFILE : medeleg:%b delegateM:%b",
	       { rg_medeleg_u1, 1'd0, rg_medeleg_m2, 2'd0, rg_medeleg_l10 },
	       rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d669 ||
	       rg_medeleg_u1_56_CONCAT_0_CONCAT_rg_medeleg_m2_ETC___d673);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d659 ||
	   TASK_testplusargs___d660 && TASK_testplusargs___d661))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d675 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d676 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d677 = $test$plusargs("l2");
	  #0;
	end
    TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d683 =
	(TASK_testplusargs___d675 ||
	 TASK_testplusargs___d676 && TASK_testplusargs___d677) &&
	rg_prv == 2'd3;
    TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d685 =
	(TASK_testplusargs___d675 ||
	 TASK_testplusargs___d676 && TASK_testplusargs___d677) &&
	rg_prv != 2'd3;
    TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d692 =
	(TASK_testplusargs___d675 ||
	 TASK_testplusargs___d676 && TASK_testplusargs___d677) &&
	NOT_rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_ETC___d691;
    TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d695 =
	(TASK_testplusargs___d675 ||
	 TASK_testplusargs___d676 && TASK_testplusargs___d677) &&
	rg_mideleg_39_SRL_upd_on_trap_cause_BITS_4_TO__ETC___d694;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  v__h14354 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d675 ||
	   TASK_testplusargs___d676 && TASK_testplusargs___d677))
	$write("[%10d", v__h14354, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d675 ||
	   TASK_testplusargs___d676 && TASK_testplusargs___d677))
	$write("CSRFILE : rg_prv: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d683)
	$write("Machine");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d685)
	$write("User");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d675 ||
	   TASK_testplusargs___d676 && TASK_testplusargs___d677))
	$write(" prv: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d692)
	$write("Machine");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  TASK_testplusargs_75_OR_TASK_testplusargs_76_A_ETC___d695)
	$write("User");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d675 ||
	   TASK_testplusargs___d676 && TASK_testplusargs___d677))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d696 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d697 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  TASK_testplusargs___d698 = $test$plusargs("l2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap)
	begin
	  v__h14564 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d696 ||
	   TASK_testplusargs___d697 && TASK_testplusargs___d698))
	$write("[%10d", v__h14564, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d696 ||
	   TASK_testplusargs___d697 && TASK_testplusargs___d698))
	$write("CSRFILE : rg_mtvec:%h rg_mode:%b", rg_mtvec, rg_mode);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_upd_on_trap &&
	  (TASK_testplusargs___d696 ||
	   TASK_testplusargs___d697 && TASK_testplusargs___d698))
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkcsrfile

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:10 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// system_instruction             O   129
// RDY_system_instruction         O     1 const
// mv_csr_decode                  O   152
// RDY_mv_csr_decode              O     1 const
// take_trap                      O    64
// RDY_take_trap                  O     1 const
// RDY_clint_msip                 O     1 const
// RDY_clint_mtip                 O     1 const
// RDY_clint_mtime                O     1 const
// RDY_incr_minstret              O     1 const
// RDY_ext_interrupt              O     1 const
// mv_csr_misa_c                  O     1 reg
// RDY_mv_csr_misa_c              O     1 const
// mv_interrupt                   O     1
// mv_curr_priv                   O     2
// RDY_mv_curr_priv               O     1 const
// csr_mstatus                    O    64
// RDY_csr_mstatus                O     1 const
// mv_pmp_cfg                     O    32 reg
// RDY_mv_pmp_cfg                 O     1 const
// mv_pmp_addr                    O   120 reg
// RDY_mv_pmp_addr                O     1 const
// mv_trigger_data1               O    44
// RDY_mv_trigger_data1           O     1 const
// mv_trigger_data2               O   128 reg
// RDY_mv_trigger_data2           O     1 const
// mv_trigger_enable              O     2
// RDY_mv_trigger_enable          O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// system_instruction_csr_address  I    12
// system_instruction_op1         I    64
// system_instruction_funct3      I     3
// system_instruction_lpc         I     2
// take_trap_type_cause           I     6
// take_trap_pc                   I    64
// take_trap_badaddr              I    64
// clint_msip_intrpt              I     1 reg
// clint_mtip_intrpt              I     1 reg
// clint_mtime_c_mtime            I    64 reg
// ext_interrupt_ex_i             I     1 reg
// EN_clint_msip                  I     1
// EN_clint_mtip                  I     1
// EN_clint_mtime                 I     1
// EN_incr_minstret               I     1
// EN_ext_interrupt               I     1
// EN_system_instruction          I     1
// EN_take_trap                   I     1
//
// Combinational paths from inputs to outputs:
//   (system_instruction_csr_address,
//    system_instruction_funct3,
//    EN_system_instruction) -> system_instruction
//   (take_trap_type_cause, EN_take_trap) -> take_trap
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkcsr(CLK,
	     RST_N,

	     system_instruction_csr_address,
	     system_instruction_op1,
	     system_instruction_funct3,
	     system_instruction_lpc,
	     EN_system_instruction,
	     system_instruction,
	     RDY_system_instruction,

	     mv_csr_decode,
	     RDY_mv_csr_decode,

	     take_trap_type_cause,
	     take_trap_pc,
	     take_trap_badaddr,
	     EN_take_trap,
	     take_trap,
	     RDY_take_trap,

	     clint_msip_intrpt,
	     EN_clint_msip,
	     RDY_clint_msip,

	     clint_mtip_intrpt,
	     EN_clint_mtip,
	     RDY_clint_mtip,

	     clint_mtime_c_mtime,
	     EN_clint_mtime,
	     RDY_clint_mtime,

	     EN_incr_minstret,
	     RDY_incr_minstret,

	     ext_interrupt_ex_i,
	     EN_ext_interrupt,
	     RDY_ext_interrupt,

	     mv_csr_misa_c,
	     RDY_mv_csr_misa_c,

	     mv_interrupt,

	     mv_curr_priv,
	     RDY_mv_curr_priv,

	     csr_mstatus,
	     RDY_csr_mstatus,

	     mv_pmp_cfg,
	     RDY_mv_pmp_cfg,

	     mv_pmp_addr,
	     RDY_mv_pmp_addr,

	     mv_trigger_data1,
	     RDY_mv_trigger_data1,

	     mv_trigger_data2,
	     RDY_mv_trigger_data2,

	     mv_trigger_enable,
	     RDY_mv_trigger_enable);
  input  CLK;
  input  RST_N;

  // actionvalue method system_instruction
  input  [11 : 0] system_instruction_csr_address;
  input  [63 : 0] system_instruction_op1;
  input  [2 : 0] system_instruction_funct3;
  input  [1 : 0] system_instruction_lpc;
  input  EN_system_instruction;
  output [128 : 0] system_instruction;
  output RDY_system_instruction;

  // value method mv_csr_decode
  output [151 : 0] mv_csr_decode;
  output RDY_mv_csr_decode;

  // actionvalue method take_trap
  input  [5 : 0] take_trap_type_cause;
  input  [63 : 0] take_trap_pc;
  input  [63 : 0] take_trap_badaddr;
  input  EN_take_trap;
  output [63 : 0] take_trap;
  output RDY_take_trap;

  // action method clint_msip
  input  clint_msip_intrpt;
  input  EN_clint_msip;
  output RDY_clint_msip;

  // action method clint_mtip
  input  clint_mtip_intrpt;
  input  EN_clint_mtip;
  output RDY_clint_mtip;

  // action method clint_mtime
  input  [63 : 0] clint_mtime_c_mtime;
  input  EN_clint_mtime;
  output RDY_clint_mtime;

  // action method incr_minstret
  input  EN_incr_minstret;
  output RDY_incr_minstret;

  // action method ext_interrupt
  input  ext_interrupt_ex_i;
  input  EN_ext_interrupt;
  output RDY_ext_interrupt;

  // value method mv_csr_misa_c
  output mv_csr_misa_c;
  output RDY_mv_csr_misa_c;

  // value method mv_interrupt
  output mv_interrupt;

  // value method mv_curr_priv
  output [1 : 0] mv_curr_priv;
  output RDY_mv_curr_priv;

  // value method csr_mstatus
  output [63 : 0] csr_mstatus;
  output RDY_csr_mstatus;

  // value method mv_pmp_cfg
  output [31 : 0] mv_pmp_cfg;
  output RDY_mv_pmp_cfg;

  // value method mv_pmp_addr
  output [119 : 0] mv_pmp_addr;
  output RDY_mv_pmp_addr;

  // value method mv_trigger_data1
  output [43 : 0] mv_trigger_data1;
  output RDY_mv_trigger_data1;

  // value method mv_trigger_data2
  output [127 : 0] mv_trigger_data2;
  output RDY_mv_trigger_data2;

  // value method mv_trigger_enable
  output [1 : 0] mv_trigger_enable;
  output RDY_mv_trigger_enable;

  // signals for module outputs
  wire [151 : 0] mv_csr_decode;
  wire [128 : 0] system_instruction;
  wire [127 : 0] mv_trigger_data2;
  wire [119 : 0] mv_pmp_addr;
  wire [63 : 0] csr_mstatus, take_trap;
  wire [43 : 0] mv_trigger_data1;
  wire [31 : 0] mv_pmp_cfg;
  wire [1 : 0] mv_curr_priv, mv_trigger_enable;
  wire RDY_clint_msip,
       RDY_clint_mtime,
       RDY_clint_mtip,
       RDY_csr_mstatus,
       RDY_ext_interrupt,
       RDY_incr_minstret,
       RDY_mv_csr_decode,
       RDY_mv_csr_misa_c,
       RDY_mv_curr_priv,
       RDY_mv_pmp_addr,
       RDY_mv_pmp_cfg,
       RDY_mv_trigger_data1,
       RDY_mv_trigger_data2,
       RDY_mv_trigger_enable,
       RDY_system_instruction,
       RDY_take_trap,
       mv_csr_misa_c,
       mv_interrupt;

  // ports of submodule csrfile
  reg [63 : 0] csrfile_write_csr_word;
  wire [151 : 0] csrfile_mv_csr_decode;
  wire [127 : 0] csrfile_mv_trigger_data2;
  wire [119 : 0] csrfile_mv_pmp_addr;
  wire [63 : 0] csrfile_clint_mtime_c_mtime,
		csrfile_csr_mstatus,
		csrfile_read_csr,
		csrfile_upd_on_ret,
		csrfile_upd_on_trap,
		csrfile_upd_on_trap_pc,
		csrfile_upd_on_trap_tval;
  wire [43 : 0] csrfile_mv_trigger_data1;
  wire [31 : 0] csrfile_mv_pmp_cfg;
  wire [11 : 0] csrfile_read_csr_addr, csrfile_write_csr_addr;
  wire [5 : 0] csrfile_upd_on_trap_cause;
  wire [1 : 0] csrfile_mv_curr_priv,
	       csrfile_mv_trigger_enable,
	       csrfile_upd_on_ret_prv,
	       csrfile_write_csr_lpc;
  wire csrfile_EN_clint_msip,
       csrfile_EN_clint_mtime,
       csrfile_EN_clint_mtip,
       csrfile_EN_ext_interrupt,
       csrfile_EN_incr_minstret,
       csrfile_EN_read_csr,
       csrfile_EN_upd_on_ret,
       csrfile_EN_upd_on_trap,
       csrfile_EN_write_csr,
       csrfile_clint_msip_intrpt,
       csrfile_clint_mtip_intrpt,
       csrfile_ext_interrupt_ex_i,
       csrfile_mv_csr_misa_c,
       csrfile_mv_interrupt;

  // rule scheduling signals
  wire CAN_FIRE_clint_msip,
       CAN_FIRE_clint_mtime,
       CAN_FIRE_clint_mtip,
       CAN_FIRE_ext_interrupt,
       CAN_FIRE_incr_minstret,
       CAN_FIRE_system_instruction,
       CAN_FIRE_take_trap,
       WILL_FIRE_clint_msip,
       WILL_FIRE_clint_mtime,
       WILL_FIRE_clint_mtip,
       WILL_FIRE_ext_interrupt,
       WILL_FIRE_incr_minstret,
       WILL_FIRE_system_instruction,
       WILL_FIRE_take_trap;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d1;
  reg TASK_testplusargs___d2;
  reg TASK_testplusargs___d3;
  reg [63 : 0] v__h434;
  reg TASK_testplusargs___d17;
  reg TASK_testplusargs___d18;
  reg TASK_testplusargs___d19;
  reg [63 : 0] v__h754;
  reg system_instruction_csr_address_BITS_11_TO_8_EQ_ETC___d22;
  // synopsys translate_on

  // remaining internal signals
  reg [63 : 0] y_avValue_snd_fst__h992;
  reg [21 : 0] CASE_csrfilemv_trigger_data1_BITS_21_TO_20_0__ETC__q2,
	       CASE_csrfilemv_trigger_data1_BITS_43_TO_42_0__ETC__q1;
  wire [63 : 0] writecsrdata__h932, writecsrdata__h933, x__h945;

  // actionvalue method system_instruction
  assign system_instruction =
	     { system_instruction_funct3 == 3'd0 &&
	       (system_instruction_csr_address[11:8] == 4'h0 ||
		system_instruction_csr_address[11:8] == 4'h3),
	       (system_instruction_funct3 == 3'd0) ?
		 { y_avValue_snd_fst__h992, 64'd0 } :
		 { 64'd0, csrfile_read_csr } } ;
  assign RDY_system_instruction = 1'd1 ;
  assign CAN_FIRE_system_instruction = 1'd1 ;
  assign WILL_FIRE_system_instruction = EN_system_instruction ;

  // value method mv_csr_decode
  assign mv_csr_decode =
	     { (csrfile_mv_csr_decode[151:150] == 2'd3) ?
		 csrfile_mv_csr_decode[151:150] :
		 2'd0,
	       csrfile_mv_csr_decode[149:0] } ;
  assign RDY_mv_csr_decode = 1'd1 ;

  // actionvalue method take_trap
  assign take_trap = csrfile_upd_on_trap ;
  assign RDY_take_trap = 1'd1 ;
  assign CAN_FIRE_take_trap = 1'd1 ;
  assign WILL_FIRE_take_trap = EN_take_trap ;

  // action method clint_msip
  assign RDY_clint_msip = 1'd1 ;
  assign CAN_FIRE_clint_msip = 1'd1 ;
  assign WILL_FIRE_clint_msip = EN_clint_msip ;

  // action method clint_mtip
  assign RDY_clint_mtip = 1'd1 ;
  assign CAN_FIRE_clint_mtip = 1'd1 ;
  assign WILL_FIRE_clint_mtip = EN_clint_mtip ;

  // action method clint_mtime
  assign RDY_clint_mtime = 1'd1 ;
  assign CAN_FIRE_clint_mtime = 1'd1 ;
  assign WILL_FIRE_clint_mtime = EN_clint_mtime ;

  // action method incr_minstret
  assign RDY_incr_minstret = 1'd1 ;
  assign CAN_FIRE_incr_minstret = 1'd1 ;
  assign WILL_FIRE_incr_minstret = EN_incr_minstret ;

  // action method ext_interrupt
  assign RDY_ext_interrupt = 1'd1 ;
  assign CAN_FIRE_ext_interrupt = 1'd1 ;
  assign WILL_FIRE_ext_interrupt = EN_ext_interrupt ;

  // value method mv_csr_misa_c
  assign mv_csr_misa_c = csrfile_mv_csr_misa_c ;
  assign RDY_mv_csr_misa_c = 1'd1 ;

  // value method mv_interrupt
  assign mv_interrupt = csrfile_mv_interrupt ;

  // value method mv_curr_priv
  assign mv_curr_priv = csrfile_mv_curr_priv ;
  assign RDY_mv_curr_priv = 1'd1 ;

  // value method csr_mstatus
  assign csr_mstatus = csrfile_csr_mstatus ;
  assign RDY_csr_mstatus = 1'd1 ;

  // value method mv_pmp_cfg
  assign mv_pmp_cfg = csrfile_mv_pmp_cfg ;
  assign RDY_mv_pmp_cfg = 1'd1 ;

  // value method mv_pmp_addr
  assign mv_pmp_addr = csrfile_mv_pmp_addr ;
  assign RDY_mv_pmp_addr = 1'd1 ;

  // value method mv_trigger_data1
  assign mv_trigger_data1 =
	     { CASE_csrfilemv_trigger_data1_BITS_43_TO_42_0__ETC__q1,
	       CASE_csrfilemv_trigger_data1_BITS_21_TO_20_0__ETC__q2 } ;
  assign RDY_mv_trigger_data1 = 1'd1 ;

  // value method mv_trigger_data2
  assign mv_trigger_data2 = csrfile_mv_trigger_data2 ;
  assign RDY_mv_trigger_data2 = 1'd1 ;

  // value method mv_trigger_enable
  assign mv_trigger_enable = csrfile_mv_trigger_enable ;
  assign RDY_mv_trigger_enable = 1'd1 ;

  // submodule csrfile
  mkcsrfile csrfile(.CLK(CLK),
		    .RST_N(RST_N),
		    .clint_msip_intrpt(csrfile_clint_msip_intrpt),
		    .clint_mtime_c_mtime(csrfile_clint_mtime_c_mtime),
		    .clint_mtip_intrpt(csrfile_clint_mtip_intrpt),
		    .ext_interrupt_ex_i(csrfile_ext_interrupt_ex_i),
		    .read_csr_addr(csrfile_read_csr_addr),
		    .upd_on_ret_prv(csrfile_upd_on_ret_prv),
		    .upd_on_trap_cause(csrfile_upd_on_trap_cause),
		    .upd_on_trap_pc(csrfile_upd_on_trap_pc),
		    .upd_on_trap_tval(csrfile_upd_on_trap_tval),
		    .write_csr_addr(csrfile_write_csr_addr),
		    .write_csr_lpc(csrfile_write_csr_lpc),
		    .write_csr_word(csrfile_write_csr_word),
		    .EN_read_csr(csrfile_EN_read_csr),
		    .EN_write_csr(csrfile_EN_write_csr),
		    .EN_upd_on_ret(csrfile_EN_upd_on_ret),
		    .EN_upd_on_trap(csrfile_EN_upd_on_trap),
		    .EN_incr_minstret(csrfile_EN_incr_minstret),
		    .EN_clint_msip(csrfile_EN_clint_msip),
		    .EN_clint_mtip(csrfile_EN_clint_mtip),
		    .EN_clint_mtime(csrfile_EN_clint_mtime),
		    .EN_ext_interrupt(csrfile_EN_ext_interrupt),
		    .read_csr(csrfile_read_csr),
		    .RDY_read_csr(),
		    .RDY_write_csr(),
		    .upd_on_ret(csrfile_upd_on_ret),
		    .RDY_upd_on_ret(),
		    .upd_on_trap(csrfile_upd_on_trap),
		    .RDY_upd_on_trap(),
		    .RDY_incr_minstret(),
		    .mv_csr_decode(csrfile_mv_csr_decode),
		    .RDY_mv_csr_decode(),
		    .mv_csr_misa_c(csrfile_mv_csr_misa_c),
		    .RDY_mv_csr_misa_c(),
		    .mv_curr_priv(csrfile_mv_curr_priv),
		    .RDY_mv_curr_priv(),
		    .csr_mstatus(csrfile_csr_mstatus),
		    .RDY_csr_mstatus(),
		    .RDY_clint_msip(),
		    .RDY_clint_mtip(),
		    .RDY_clint_mtime(),
		    .RDY_ext_interrupt(),
		    .mv_interrupt(csrfile_mv_interrupt),
		    .mv_pmp_cfg(csrfile_mv_pmp_cfg),
		    .RDY_mv_pmp_cfg(),
		    .mv_pmp_addr(csrfile_mv_pmp_addr),
		    .RDY_mv_pmp_addr(),
		    .mv_trigger_data1(csrfile_mv_trigger_data1),
		    .RDY_mv_trigger_data1(),
		    .mv_trigger_data2(csrfile_mv_trigger_data2),
		    .RDY_mv_trigger_data2(),
		    .mv_trigger_enable(csrfile_mv_trigger_enable),
		    .RDY_mv_trigger_enable());

  // submodule csrfile
  assign csrfile_clint_msip_intrpt = clint_msip_intrpt ;
  assign csrfile_clint_mtime_c_mtime = clint_mtime_c_mtime ;
  assign csrfile_clint_mtip_intrpt = clint_mtip_intrpt ;
  assign csrfile_ext_interrupt_ex_i = ext_interrupt_ex_i ;
  assign csrfile_read_csr_addr = system_instruction_csr_address ;
  assign csrfile_upd_on_ret_prv =
	     (system_instruction_csr_address[9:8] == 2'd3) ?
	       system_instruction_csr_address[9:8] :
	       2'd0 ;
  assign csrfile_upd_on_trap_cause = take_trap_type_cause ;
  assign csrfile_upd_on_trap_pc = take_trap_pc ;
  assign csrfile_upd_on_trap_tval = take_trap_badaddr ;
  assign csrfile_write_csr_addr = system_instruction_csr_address ;
  assign csrfile_write_csr_lpc = system_instruction_lpc ;
  always@(system_instruction_funct3 or
	  writecsrdata__h933 or system_instruction_op1 or writecsrdata__h932)
  begin
    case (system_instruction_funct3[1:0])
      2'd1: csrfile_write_csr_word = system_instruction_op1;
      2'd2: csrfile_write_csr_word = writecsrdata__h932;
      default: csrfile_write_csr_word = writecsrdata__h933;
    endcase
  end
  assign csrfile_EN_read_csr = EN_system_instruction ;
  assign csrfile_EN_write_csr =
	     EN_system_instruction && system_instruction_funct3 != 3'd0 ;
  assign csrfile_EN_upd_on_ret =
	     EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	     (system_instruction_csr_address[11:8] == 4'h0 ||
	      system_instruction_csr_address[11:8] == 4'h3) ;
  assign csrfile_EN_upd_on_trap = EN_take_trap ;
  assign csrfile_EN_incr_minstret = EN_incr_minstret ;
  assign csrfile_EN_clint_msip = EN_clint_msip ;
  assign csrfile_EN_clint_mtip = EN_clint_mtip ;
  assign csrfile_EN_clint_mtime = EN_clint_mtime ;
  assign csrfile_EN_ext_interrupt = EN_ext_interrupt ;

  // remaining internal signals
  assign writecsrdata__h932 = system_instruction_op1 | csrfile_read_csr ;
  assign writecsrdata__h933 = x__h945 & csrfile_read_csr ;
  assign x__h945 = ~system_instruction_op1 ;
  always@(csrfile_mv_trigger_data1)
  begin
    case (csrfile_mv_trigger_data1[43:42])
      2'd0, 2'd1, 2'd2:
	  CASE_csrfilemv_trigger_data1_BITS_43_TO_42_0__ETC__q1 =
	      csrfile_mv_trigger_data1[43:22];
      2'd3:
	  CASE_csrfilemv_trigger_data1_BITS_43_TO_42_0__ETC__q1 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(csrfile_mv_trigger_data1)
  begin
    case (csrfile_mv_trigger_data1[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_csrfilemv_trigger_data1_BITS_21_TO_20_0__ETC__q2 =
	      csrfile_mv_trigger_data1[21:0];
      2'd3:
	  CASE_csrfilemv_trigger_data1_BITS_21_TO_20_0__ETC__q2 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(system_instruction_csr_address or csrfile_upd_on_ret)
  begin
    case (system_instruction_csr_address[11:8])
      4'h0, 4'h3: y_avValue_snd_fst__h992 = csrfile_upd_on_ret;
      default: y_avValue_snd_fst__h992 = 64'd0;
    endcase
  end

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction)
	begin
	  TASK_testplusargs___d1 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction)
	begin
	  TASK_testplusargs___d2 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction)
	begin
	  TASK_testplusargs___d3 = $test$plusargs("l2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction)
	begin
	  v__h434 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction &&
	  (TASK_testplusargs___d1 ||
	   TASK_testplusargs___d2 && TASK_testplusargs___d3))
	$write("[%10d", v__h434, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction &&
	  (TASK_testplusargs___d1 ||
	   TASK_testplusargs___d2 && TASK_testplusargs___d3))
	$write("CSR : Operation csr: %h op1: %h, funct3: %b csr_read: %h",
	       system_instruction_csr_address,
	       system_instruction_op1,
	       system_instruction_funct3,
	       csrfile_read_csr);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction &&
	  (TASK_testplusargs___d1 ||
	   TASK_testplusargs___d2 && TASK_testplusargs___d3))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  (system_instruction_csr_address[11:8] == 4'h0 ||
	   system_instruction_csr_address[11:8] == 4'h3))
	begin
	  TASK_testplusargs___d17 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  (system_instruction_csr_address[11:8] == 4'h0 ||
	   system_instruction_csr_address[11:8] == 4'h3))
	begin
	  TASK_testplusargs___d18 = $test$plusargs("mcsr");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  (system_instruction_csr_address[11:8] == 4'h0 ||
	   system_instruction_csr_address[11:8] == 4'h3))
	begin
	  TASK_testplusargs___d19 = $test$plusargs("l1");
	  #0;
	end
    system_instruction_csr_address_BITS_11_TO_8_EQ_ETC___d22 =
	(system_instruction_csr_address[11:8] == 4'h0 ||
	 system_instruction_csr_address[11:8] == 4'h3) &&
	(TASK_testplusargs___d17 ||
	 TASK_testplusargs___d18 && TASK_testplusargs___d19);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  (system_instruction_csr_address[11:8] == 4'h0 ||
	   system_instruction_csr_address[11:8] == 4'h3))
	begin
	  v__h754 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  system_instruction_csr_address_BITS_11_TO_8_EQ_ETC___d22)
	$write("[%10d", v__h754, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  system_instruction_csr_address_BITS_11_TO_8_EQ_ETC___d22)
	$write("CSR : RET Function: %h", system_instruction_csr_address);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_system_instruction && system_instruction_funct3 == 3'd0 &&
	  system_instruction_csr_address_BITS_11_TO_8_EQ_ETC___d22)
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkcsr

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:18 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// master_d_awvalid               O     1 reg
// master_d_awaddr                O    32 reg
// master_d_awprot                O     3 reg
// master_d_awsize                O     2 reg
// master_d_wvalid                O     1 reg
// master_d_wdata                 O    64 reg
// master_d_wstrb                 O     8 reg
// master_d_bready                O     1 reg
// master_d_arvalid               O     1 reg
// master_d_araddr                O    32 reg
// master_d_arprot                O     3 reg
// master_d_arsize                O     2 reg
// master_d_rready                O     1 reg
// master_i_awvalid               O     1 reg
// master_i_awaddr                O    32 reg
// master_i_awprot                O     3 reg
// master_i_awsize                O     2 reg
// master_i_wvalid                O     1 reg
// master_i_wdata                 O    64 reg
// master_i_wstrb                 O     8 reg
// master_i_bready                O     1 reg
// master_i_arvalid               O     1 reg
// master_i_araddr                O    32 reg
// master_i_arprot                O     3 reg
// master_i_arsize                O     2 reg
// master_i_rready                O     1 reg
// RDY_sb_clint_msip_put          O     1 const
// RDY_sb_clint_mtip_put          O     1 const
// RDY_sb_clint_mtime_put         O     1 const
// RDY_sb_ext_interrupt_put       O     1 const
// io_dump_get                    O   167
// RDY_io_dump_get                O     1 reg
// resetpc                        I    64
// CLK                            I     1 clock
// RST_N                          I     1 reset
// master_d_m_awready_awready     I     1
// master_d_m_wready_wready       I     1
// master_d_m_bvalid_bvalid       I     1
// master_d_m_bvalid_bresp        I     2 reg
// master_d_m_arready_arready     I     1
// master_d_m_rvalid_rvalid       I     1
// master_d_m_rvalid_rresp        I     2 reg
// master_d_m_rvalid_rdata        I    64 reg
// master_i_m_awready_awready     I     1
// master_i_m_wready_wready       I     1
// master_i_m_bvalid_bvalid       I     1
// master_i_m_bvalid_bresp        I     2 reg
// master_i_m_arready_arready     I     1
// master_i_m_rvalid_rvalid       I     1
// master_i_m_rvalid_rresp        I     2 reg
// master_i_m_rvalid_rdata        I    64 reg
// sb_clint_msip_put              I     1 reg
// sb_clint_mtip_put              I     1 reg
// sb_clint_mtime_put             I    64 reg
// sb_ext_interrupt_put           I     1 reg
// EN_sb_clint_msip_put           I     1
// EN_sb_clint_mtip_put           I     1
// EN_sb_clint_mtime_put          I     1
// EN_sb_ext_interrupt_put        I     1
// EN_io_dump_get                 I     1
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkeclass_axi4lite(resetpc,
			 CLK,
			 RST_N,

			 master_d_awvalid,

			 master_d_awaddr,

			 master_d_awprot,

			 master_d_awsize,

			 master_d_m_awready_awready,

			 master_d_wvalid,

			 master_d_wdata,

			 master_d_wstrb,

			 master_d_m_wready_wready,

			 master_d_m_bvalid_bvalid,
			 master_d_m_bvalid_bresp,

			 master_d_bready,

			 master_d_arvalid,

			 master_d_araddr,

			 master_d_arprot,

			 master_d_arsize,

			 master_d_m_arready_arready,

			 master_d_m_rvalid_rvalid,
			 master_d_m_rvalid_rresp,
			 master_d_m_rvalid_rdata,

			 master_d_rready,

			 master_i_awvalid,

			 master_i_awaddr,

			 master_i_awprot,

			 master_i_awsize,

			 master_i_m_awready_awready,

			 master_i_wvalid,

			 master_i_wdata,

			 master_i_wstrb,

			 master_i_m_wready_wready,

			 master_i_m_bvalid_bvalid,
			 master_i_m_bvalid_bresp,

			 master_i_bready,

			 master_i_arvalid,

			 master_i_araddr,

			 master_i_arprot,

			 master_i_arsize,

			 master_i_m_arready_arready,

			 master_i_m_rvalid_rvalid,
			 master_i_m_rvalid_rresp,
			 master_i_m_rvalid_rdata,

			 master_i_rready,

			 sb_clint_msip_put,
			 EN_sb_clint_msip_put,
			 RDY_sb_clint_msip_put,

			 sb_clint_mtip_put,
			 EN_sb_clint_mtip_put,
			 RDY_sb_clint_mtip_put,

			 sb_clint_mtime_put,
			 EN_sb_clint_mtime_put,
			 RDY_sb_clint_mtime_put,

			 sb_ext_interrupt_put,
			 EN_sb_ext_interrupt_put,
			 RDY_sb_ext_interrupt_put,

			 EN_io_dump_get,
			 io_dump_get,
			 RDY_io_dump_get);
  input  [63 : 0] resetpc;
  input  CLK;
  input  RST_N;

  // value method master_d_m_awvalid
  output master_d_awvalid;

  // value method master_d_m_awaddr
  output [31 : 0] master_d_awaddr;

  // value method master_d_m_awuser

  // value method master_d_m_awprot
  output [2 : 0] master_d_awprot;

  // value method master_d_m_awsize
  output [1 : 0] master_d_awsize;

  // action method master_d_m_awready
  input  master_d_m_awready_awready;

  // value method master_d_m_wvalid
  output master_d_wvalid;

  // value method master_d_m_wdata
  output [63 : 0] master_d_wdata;

  // value method master_d_m_wstrb
  output [7 : 0] master_d_wstrb;

  // action method master_d_m_wready
  input  master_d_m_wready_wready;

  // action method master_d_m_bvalid
  input  master_d_m_bvalid_bvalid;
  input  [1 : 0] master_d_m_bvalid_bresp;

  // value method master_d_m_bready
  output master_d_bready;

  // value method master_d_m_arvalid
  output master_d_arvalid;

  // value method master_d_m_araddr
  output [31 : 0] master_d_araddr;

  // value method master_d_m_aruser

  // value method master_d_m_arprot
  output [2 : 0] master_d_arprot;

  // value method master_d_m_arsize
  output [1 : 0] master_d_arsize;

  // action method master_d_m_arready
  input  master_d_m_arready_arready;

  // action method master_d_m_rvalid
  input  master_d_m_rvalid_rvalid;
  input  [1 : 0] master_d_m_rvalid_rresp;
  input  [63 : 0] master_d_m_rvalid_rdata;

  // value method master_d_m_rready
  output master_d_rready;

  // value method master_i_m_awvalid
  output master_i_awvalid;

  // value method master_i_m_awaddr
  output [31 : 0] master_i_awaddr;

  // value method master_i_m_awuser

  // value method master_i_m_awprot
  output [2 : 0] master_i_awprot;

  // value method master_i_m_awsize
  output [1 : 0] master_i_awsize;

  // action method master_i_m_awready
  input  master_i_m_awready_awready;

  // value method master_i_m_wvalid
  output master_i_wvalid;

  // value method master_i_m_wdata
  output [63 : 0] master_i_wdata;

  // value method master_i_m_wstrb
  output [7 : 0] master_i_wstrb;

  // action method master_i_m_wready
  input  master_i_m_wready_wready;

  // action method master_i_m_bvalid
  input  master_i_m_bvalid_bvalid;
  input  [1 : 0] master_i_m_bvalid_bresp;

  // value method master_i_m_bready
  output master_i_bready;

  // value method master_i_m_arvalid
  output master_i_arvalid;

  // value method master_i_m_araddr
  output [31 : 0] master_i_araddr;

  // value method master_i_m_aruser

  // value method master_i_m_arprot
  output [2 : 0] master_i_arprot;

  // value method master_i_m_arsize
  output [1 : 0] master_i_arsize;

  // action method master_i_m_arready
  input  master_i_m_arready_arready;

  // action method master_i_m_rvalid
  input  master_i_m_rvalid_rvalid;
  input  [1 : 0] master_i_m_rvalid_rresp;
  input  [63 : 0] master_i_m_rvalid_rdata;

  // value method master_i_m_rready
  output master_i_rready;

  // action method sb_clint_msip_put
  input  sb_clint_msip_put;
  input  EN_sb_clint_msip_put;
  output RDY_sb_clint_msip_put;

  // action method sb_clint_mtip_put
  input  sb_clint_mtip_put;
  input  EN_sb_clint_mtip_put;
  output RDY_sb_clint_mtip_put;

  // action method sb_clint_mtime_put
  input  [63 : 0] sb_clint_mtime_put;
  input  EN_sb_clint_mtime_put;
  output RDY_sb_clint_mtime_put;

  // action method sb_ext_interrupt_put
  input  sb_ext_interrupt_put;
  input  EN_sb_ext_interrupt_put;
  output RDY_sb_ext_interrupt_put;

  // actionvalue method io_dump_get
  input  EN_io_dump_get;
  output [166 : 0] io_dump_get;
  output RDY_io_dump_get;

  // signals for module outputs
  wire [166 : 0] io_dump_get;
  wire [63 : 0] master_d_wdata, master_i_wdata;
  wire [31 : 0] master_d_araddr,
		master_d_awaddr,
		master_i_araddr,
		master_i_awaddr;
  wire [7 : 0] master_d_wstrb, master_i_wstrb;
  wire [2 : 0] master_d_arprot,
	       master_d_awprot,
	       master_i_arprot,
	       master_i_awprot;
  wire [1 : 0] master_d_arsize,
	       master_d_awsize,
	       master_i_arsize,
	       master_i_awsize;
  wire RDY_io_dump_get,
       RDY_sb_clint_msip_put,
       RDY_sb_clint_mtime_put,
       RDY_sb_clint_mtip_put,
       RDY_sb_ext_interrupt_put,
       master_d_arvalid,
       master_d_awvalid,
       master_d_bready,
       master_d_rready,
       master_d_wvalid,
       master_i_arvalid,
       master_i_awvalid,
       master_i_bready,
       master_i_rready,
       master_i_wvalid;

  // register rg_wEpoch
  reg rg_wEpoch;
  wire rg_wEpoch_D_IN, rg_wEpoch_EN;

  // ports of submodule fetch_xactor_f_rd_addr
  wire [36 : 0] fetch_xactor_f_rd_addr_D_IN, fetch_xactor_f_rd_addr_D_OUT;
  wire fetch_xactor_f_rd_addr_CLR,
       fetch_xactor_f_rd_addr_DEQ,
       fetch_xactor_f_rd_addr_EMPTY_N,
       fetch_xactor_f_rd_addr_ENQ,
       fetch_xactor_f_rd_addr_FULL_N;

  // ports of submodule fetch_xactor_f_rd_data
  wire [65 : 0] fetch_xactor_f_rd_data_D_IN, fetch_xactor_f_rd_data_D_OUT;
  wire fetch_xactor_f_rd_data_CLR,
       fetch_xactor_f_rd_data_DEQ,
       fetch_xactor_f_rd_data_EMPTY_N,
       fetch_xactor_f_rd_data_ENQ,
       fetch_xactor_f_rd_data_FULL_N;

  // ports of submodule fetch_xactor_f_wr_addr
  wire [36 : 0] fetch_xactor_f_wr_addr_D_IN, fetch_xactor_f_wr_addr_D_OUT;
  wire fetch_xactor_f_wr_addr_CLR,
       fetch_xactor_f_wr_addr_DEQ,
       fetch_xactor_f_wr_addr_EMPTY_N,
       fetch_xactor_f_wr_addr_ENQ;

  // ports of submodule fetch_xactor_f_wr_data
  wire [71 : 0] fetch_xactor_f_wr_data_D_IN, fetch_xactor_f_wr_data_D_OUT;
  wire fetch_xactor_f_wr_data_CLR,
       fetch_xactor_f_wr_data_DEQ,
       fetch_xactor_f_wr_data_EMPTY_N,
       fetch_xactor_f_wr_data_ENQ;

  // ports of submodule fetch_xactor_f_wr_resp
  wire [1 : 0] fetch_xactor_f_wr_resp_D_IN;
  wire fetch_xactor_f_wr_resp_CLR,
       fetch_xactor_f_wr_resp_DEQ,
       fetch_xactor_f_wr_resp_ENQ,
       fetch_xactor_f_wr_resp_FULL_N;

  // ports of submodule ff_atomic_state
  wire [63 : 0] ff_atomic_state_D_IN, ff_atomic_state_D_OUT;
  wire ff_atomic_state_CLR,
       ff_atomic_state_DEQ,
       ff_atomic_state_EMPTY_N,
       ff_atomic_state_ENQ,
       ff_atomic_state_FULL_N;

  // ports of submodule ff_inst_access_fault
  wire ff_inst_access_fault_CLR,
       ff_inst_access_fault_DEQ,
       ff_inst_access_fault_D_IN,
       ff_inst_access_fault_D_OUT,
       ff_inst_access_fault_EMPTY_N,
       ff_inst_access_fault_ENQ,
       ff_inst_access_fault_FULL_N;

  // ports of submodule ff_inst_request
  wire [65 : 0] ff_inst_request_D_IN, ff_inst_request_D_OUT;
  wire ff_inst_request_CLR,
       ff_inst_request_DEQ,
       ff_inst_request_EMPTY_N,
       ff_inst_request_ENQ,
       ff_inst_request_FULL_N;

  // ports of submodule ff_mem_access_fault
  wire ff_mem_access_fault_CLR,
       ff_mem_access_fault_DEQ,
       ff_mem_access_fault_D_IN,
       ff_mem_access_fault_ENQ;

  // ports of submodule ff_mem_request
  wire [138 : 0] ff_mem_request_D_IN, ff_mem_request_D_OUT;
  wire ff_mem_request_CLR,
       ff_mem_request_DEQ,
       ff_mem_request_EMPTY_N,
       ff_mem_request_ENQ,
       ff_mem_request_FULL_N;

  // ports of submodule memory_xactor_f_rd_addr
  wire [36 : 0] memory_xactor_f_rd_addr_D_IN, memory_xactor_f_rd_addr_D_OUT;
  wire memory_xactor_f_rd_addr_CLR,
       memory_xactor_f_rd_addr_DEQ,
       memory_xactor_f_rd_addr_EMPTY_N,
       memory_xactor_f_rd_addr_ENQ,
       memory_xactor_f_rd_addr_FULL_N;

  // ports of submodule memory_xactor_f_rd_data
  wire [65 : 0] memory_xactor_f_rd_data_D_IN, memory_xactor_f_rd_data_D_OUT;
  wire memory_xactor_f_rd_data_CLR,
       memory_xactor_f_rd_data_DEQ,
       memory_xactor_f_rd_data_EMPTY_N,
       memory_xactor_f_rd_data_ENQ,
       memory_xactor_f_rd_data_FULL_N;

  // ports of submodule memory_xactor_f_wr_addr
  wire [36 : 0] memory_xactor_f_wr_addr_D_IN, memory_xactor_f_wr_addr_D_OUT;
  wire memory_xactor_f_wr_addr_CLR,
       memory_xactor_f_wr_addr_DEQ,
       memory_xactor_f_wr_addr_EMPTY_N,
       memory_xactor_f_wr_addr_ENQ,
       memory_xactor_f_wr_addr_FULL_N;

  // ports of submodule memory_xactor_f_wr_data
  wire [71 : 0] memory_xactor_f_wr_data_D_IN, memory_xactor_f_wr_data_D_OUT;
  wire memory_xactor_f_wr_data_CLR,
       memory_xactor_f_wr_data_DEQ,
       memory_xactor_f_wr_data_EMPTY_N,
       memory_xactor_f_wr_data_ENQ,
       memory_xactor_f_wr_data_FULL_N;

  // ports of submodule memory_xactor_f_wr_resp
  wire [1 : 0] memory_xactor_f_wr_resp_D_IN, memory_xactor_f_wr_resp_D_OUT;
  wire memory_xactor_f_wr_resp_CLR,
       memory_xactor_f_wr_resp_DEQ,
       memory_xactor_f_wr_resp_EMPTY_N,
       memory_xactor_f_wr_resp_ENQ,
       memory_xactor_f_wr_resp_FULL_N;

  // ports of submodule riscv
  reg [65 : 0] riscv_memory_response_put;
  wire [166 : 0] riscv_dump_get;
  wire [138 : 0] riscv_memory_request_get;
  wire [119 : 0] riscv_mv_pmp_addr;
  wire [65 : 0] riscv_inst_request_get;
  wire [63 : 0] riscv_clint_mtime_c_mtime;
  wire [34 : 0] riscv_inst_response_put;
  wire [31 : 0] riscv_mv_pmp_cfg;
  wire [1 : 0] riscv_mv_curr_priv;
  wire riscv_EN_clint_msip,
       riscv_EN_clint_mtime,
       riscv_EN_clint_mtip,
       riscv_EN_dump_get,
       riscv_EN_ext_interrupt,
       riscv_EN_inst_request_get,
       riscv_EN_inst_response_put,
       riscv_EN_memory_request_get,
       riscv_EN_memory_response_put,
       riscv_RDY_dump_get,
       riscv_RDY_inst_request_get,
       riscv_RDY_inst_response_put,
       riscv_RDY_memory_request_get,
       riscv_clint_msip_intrpt,
       riscv_clint_mtip_intrpt,
       riscv_ext_interrupt_intrpt,
       riscv_mv_trap;

  // rule scheduling signals
  wire CAN_FIRE_RL_handle_atomic_readresponse,
       CAN_FIRE_RL_handle_atomic_writeresponse,
       CAN_FIRE_RL_handle_fetch_request,
       CAN_FIRE_RL_handle_fetch_response,
       CAN_FIRE_RL_handle_inst_access_fault,
       CAN_FIRE_RL_handle_memoryRead_response,
       CAN_FIRE_RL_handle_memoryWrite_response,
       CAN_FIRE_RL_handle_memory_request,
       CAN_FIRE_RL_update_epochs,
       CAN_FIRE_io_dump_get,
       CAN_FIRE_master_d_m_arready,
       CAN_FIRE_master_d_m_awready,
       CAN_FIRE_master_d_m_bvalid,
       CAN_FIRE_master_d_m_rvalid,
       CAN_FIRE_master_d_m_wready,
       CAN_FIRE_master_i_m_arready,
       CAN_FIRE_master_i_m_awready,
       CAN_FIRE_master_i_m_bvalid,
       CAN_FIRE_master_i_m_rvalid,
       CAN_FIRE_master_i_m_wready,
       CAN_FIRE_sb_clint_msip_put,
       CAN_FIRE_sb_clint_mtime_put,
       CAN_FIRE_sb_clint_mtip_put,
       CAN_FIRE_sb_ext_interrupt_put,
       WILL_FIRE_RL_handle_atomic_readresponse,
       WILL_FIRE_RL_handle_atomic_writeresponse,
       WILL_FIRE_RL_handle_fetch_request,
       WILL_FIRE_RL_handle_fetch_response,
       WILL_FIRE_RL_handle_inst_access_fault,
       WILL_FIRE_RL_handle_memoryRead_response,
       WILL_FIRE_RL_handle_memoryWrite_response,
       WILL_FIRE_RL_handle_memory_request,
       WILL_FIRE_RL_update_epochs,
       WILL_FIRE_io_dump_get,
       WILL_FIRE_master_d_m_arready,
       WILL_FIRE_master_d_m_awready,
       WILL_FIRE_master_d_m_bvalid,
       WILL_FIRE_master_d_m_rvalid,
       WILL_FIRE_master_d_m_wready,
       WILL_FIRE_master_i_m_arready,
       WILL_FIRE_master_i_m_awready,
       WILL_FIRE_master_i_m_bvalid,
       WILL_FIRE_master_i_m_rvalid,
       WILL_FIRE_master_i_m_wready,
       WILL_FIRE_sb_clint_msip_put,
       WILL_FIRE_sb_clint_mtime_put,
       WILL_FIRE_sb_clint_mtip_put,
       WILL_FIRE_sb_ext_interrupt_put;

  // inputs to muxes for submodule ports
  wire [71 : 0] MUX_memory_xactor_f_wr_data_enq_1__VAL_1,
		MUX_memory_xactor_f_wr_data_enq_1__VAL_2;
  wire [65 : 0] MUX_riscv_memory_response_put_1__VAL_1,
		MUX_riscv_memory_response_put_1__VAL_2,
		MUX_riscv_memory_response_put_1__VAL_3,
		MUX_riscv_memory_response_put_1__VAL_4;
  wire [36 : 0] MUX_memory_xactor_f_wr_addr_enq_1__VAL_1,
		MUX_memory_xactor_f_wr_addr_enq_1__VAL_2;
  wire [34 : 0] MUX_riscv_inst_response_put_1__VAL_1,
		MUX_riscv_inst_response_put_1__VAL_2;
  wire MUX_memory_xactor_f_wr_addr_enq_1__SEL_1,
       MUX_riscv_memory_response_put_1__SEL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d28;
  reg TASK_testplusargs___d29;
  reg TASK_testplusargs___d30;
  reg [63 : 0] v__h3195;
  reg TASK_testplusargs___d37;
  reg TASK_testplusargs___d38;
  reg TASK_testplusargs___d39;
  reg [63 : 0] v__h3370;
  reg TASK_testplusargs___d70;
  reg TASK_testplusargs___d71;
  reg TASK_testplusargs___d72;
  reg [63 : 0] v__h3802;
  reg TASK_testplusargs___d91;
  reg TASK_testplusargs___d92;
  reg TASK_testplusargs___d93;
  reg [63 : 0] v__h4000;
  reg TASK_testplusargs___d154;
  reg TASK_testplusargs___d155;
  reg TASK_testplusargs___d156;
  reg [63 : 0] v__h7409;
  reg TASK_testplusargs___d162;
  reg TASK_testplusargs___d163;
  reg TASK_testplusargs___d164;
  reg [63 : 0] v__h7569;
  reg TASK_testplusargs___d172;
  reg TASK_testplusargs___d173;
  reg TASK_testplusargs___d174;
  reg [63 : 0] v__h5179;
  reg TASK_testplusargs___d227;
  reg TASK_testplusargs___d228;
  reg TASK_testplusargs___d229;
  reg [63 : 0] v__h8304;
  reg TASK_testplusargs___d253;
  reg TASK_testplusargs___d254;
  reg TASK_testplusargs___d255;
  reg [63 : 0] v__h8610;
  reg TASK_testplusargs___d284;
  reg TASK_testplusargs___d285;
  reg TASK_testplusargs___d286;
  reg [63 : 0] v__h8793;
  reg TASK_testplusargs___d351;
  reg TASK_testplusargs___d352;
  reg TASK_testplusargs___d353;
  reg [63 : 0] v__h10105;
  reg riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159;
  reg riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167;
  reg NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177;
  reg riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33;
  reg NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42;
  reg TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d76;
  reg TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d78;
  reg TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d80;
  reg TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d85;
  reg TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d233;
  reg TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d235;
  reg TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d237;
  reg TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d242;
  reg TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d259;
  reg TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d261;
  reg TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d263;
  reg TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d268;
  reg TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d290;
  reg TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d291;
  reg TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d292;
  reg TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d293;
  reg TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d357;
  reg TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d358;
  reg TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d359;
  reg TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d360;
  // synopsys translate_on

  // remaining internal signals
  reg [63 : 0] IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220,
	       w_wdata__h5384,
	       wdata__h9103;
  reg [7 : 0] write_strobe__h4071;
  reg [1 : 0] CASE_riscvmemory_request_get_BITS_10_TO_9_0_r_ETC__q6;
  wire [63 : 0] IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d218,
		IF_ff_mem_request_first__90_BIT_8_99_THEN_0_CO_ETC___d217,
		lv_data__h3600,
		op1___1__h9539,
		op1__h9481,
		op2___1__h9540,
		op2__h9482,
		put_data__h7891,
		put_data__h8506,
		put_data__h9976,
		rdata__h7865,
		wdata___1__h9203,
		x__h3633,
		x__h5078;
  wire [31 : 0] IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC__q3,
		ff_mem_requestD_OUT_BITS_42_TO_11__q1,
		pmpreq_address__h1928,
		pmpreq_address__h4100,
		rdata865_BITS_31_TO_0__q2;
  wire [15 : 0] rdata865_BITS_15_TO_0__q5;
  wire [7 : 0] rdata865_BITS_7_TO_0__q4,
	       w_wstrb__h5385,
	       write_strobe___1__h7282,
	       write_strobe___1__h9202,
	       write_strobe__h8725;
  wire [6 : 0] fn_pmp_lookup___d119, fn_pmp_lookup___d21;
  wire [5 : 0] lv_shift__h3599, lv_shift__h7864, pmpreq_num_bytes__h4101;
  wire [2 : 0] aw_awprot__h9129;
  wire [1 : 0] IF_riscv_mv_curr_priv__6_EQ_3_7_THEN_riscv_mv__ETC___d18,
	       pmpreq_access_type__h4102;
  wire IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d317,
       IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d322,
       rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109,
       x_port1__read__h4086;

  // value method master_d_m_awvalid
  assign master_d_awvalid = memory_xactor_f_wr_addr_EMPTY_N ;

  // value method master_d_m_awaddr
  assign master_d_awaddr = memory_xactor_f_wr_addr_D_OUT[36:5] ;

  // value method master_d_m_awprot
  assign master_d_awprot = memory_xactor_f_wr_addr_D_OUT[4:2] ;

  // value method master_d_m_awsize
  assign master_d_awsize = memory_xactor_f_wr_addr_D_OUT[1:0] ;

  // action method master_d_m_awready
  assign CAN_FIRE_master_d_m_awready = 1'd1 ;
  assign WILL_FIRE_master_d_m_awready = 1'd1 ;

  // value method master_d_m_wvalid
  assign master_d_wvalid = memory_xactor_f_wr_data_EMPTY_N ;

  // value method master_d_m_wdata
  assign master_d_wdata = memory_xactor_f_wr_data_D_OUT[71:8] ;

  // value method master_d_m_wstrb
  assign master_d_wstrb = memory_xactor_f_wr_data_D_OUT[7:0] ;

  // action method master_d_m_wready
  assign CAN_FIRE_master_d_m_wready = 1'd1 ;
  assign WILL_FIRE_master_d_m_wready = 1'd1 ;

  // action method master_d_m_bvalid
  assign CAN_FIRE_master_d_m_bvalid = 1'd1 ;
  assign WILL_FIRE_master_d_m_bvalid = 1'd1 ;

  // value method master_d_m_bready
  assign master_d_bready = memory_xactor_f_wr_resp_FULL_N ;

  // value method master_d_m_arvalid
  assign master_d_arvalid = memory_xactor_f_rd_addr_EMPTY_N ;

  // value method master_d_m_araddr
  assign master_d_araddr = memory_xactor_f_rd_addr_D_OUT[36:5] ;

  // value method master_d_m_arprot
  assign master_d_arprot = memory_xactor_f_rd_addr_D_OUT[4:2] ;

  // value method master_d_m_arsize
  assign master_d_arsize = memory_xactor_f_rd_addr_D_OUT[1:0] ;

  // action method master_d_m_arready
  assign CAN_FIRE_master_d_m_arready = 1'd1 ;
  assign WILL_FIRE_master_d_m_arready = 1'd1 ;

  // action method master_d_m_rvalid
  assign CAN_FIRE_master_d_m_rvalid = 1'd1 ;
  assign WILL_FIRE_master_d_m_rvalid = 1'd1 ;

  // value method master_d_m_rready
  assign master_d_rready = memory_xactor_f_rd_data_FULL_N ;

  // value method master_i_m_awvalid
  assign master_i_awvalid = fetch_xactor_f_wr_addr_EMPTY_N ;

  // value method master_i_m_awaddr
  assign master_i_awaddr = fetch_xactor_f_wr_addr_D_OUT[36:5] ;

  // value method master_i_m_awprot
  assign master_i_awprot = fetch_xactor_f_wr_addr_D_OUT[4:2] ;

  // value method master_i_m_awsize
  assign master_i_awsize = fetch_xactor_f_wr_addr_D_OUT[1:0] ;

  // action method master_i_m_awready
  assign CAN_FIRE_master_i_m_awready = 1'd1 ;
  assign WILL_FIRE_master_i_m_awready = 1'd1 ;

  // value method master_i_m_wvalid
  assign master_i_wvalid = fetch_xactor_f_wr_data_EMPTY_N ;

  // value method master_i_m_wdata
  assign master_i_wdata = fetch_xactor_f_wr_data_D_OUT[71:8] ;

  // value method master_i_m_wstrb
  assign master_i_wstrb = fetch_xactor_f_wr_data_D_OUT[7:0] ;

  // action method master_i_m_wready
  assign CAN_FIRE_master_i_m_wready = 1'd1 ;
  assign WILL_FIRE_master_i_m_wready = 1'd1 ;

  // action method master_i_m_bvalid
  assign CAN_FIRE_master_i_m_bvalid = 1'd1 ;
  assign WILL_FIRE_master_i_m_bvalid = 1'd1 ;

  // value method master_i_m_bready
  assign master_i_bready = fetch_xactor_f_wr_resp_FULL_N ;

  // value method master_i_m_arvalid
  assign master_i_arvalid = fetch_xactor_f_rd_addr_EMPTY_N ;

  // value method master_i_m_araddr
  assign master_i_araddr = fetch_xactor_f_rd_addr_D_OUT[36:5] ;

  // value method master_i_m_arprot
  assign master_i_arprot = fetch_xactor_f_rd_addr_D_OUT[4:2] ;

  // value method master_i_m_arsize
  assign master_i_arsize = fetch_xactor_f_rd_addr_D_OUT[1:0] ;

  // action method master_i_m_arready
  assign CAN_FIRE_master_i_m_arready = 1'd1 ;
  assign WILL_FIRE_master_i_m_arready = 1'd1 ;

  // action method master_i_m_rvalid
  assign CAN_FIRE_master_i_m_rvalid = 1'd1 ;
  assign WILL_FIRE_master_i_m_rvalid = 1'd1 ;

  // value method master_i_m_rready
  assign master_i_rready = fetch_xactor_f_rd_data_FULL_N ;

  // action method sb_clint_msip_put
  assign RDY_sb_clint_msip_put = 1'd1 ;
  assign CAN_FIRE_sb_clint_msip_put = 1'd1 ;
  assign WILL_FIRE_sb_clint_msip_put = EN_sb_clint_msip_put ;

  // action method sb_clint_mtip_put
  assign RDY_sb_clint_mtip_put = 1'd1 ;
  assign CAN_FIRE_sb_clint_mtip_put = 1'd1 ;
  assign WILL_FIRE_sb_clint_mtip_put = EN_sb_clint_mtip_put ;

  // action method sb_clint_mtime_put
  assign RDY_sb_clint_mtime_put = 1'd1 ;
  assign CAN_FIRE_sb_clint_mtime_put = 1'd1 ;
  assign WILL_FIRE_sb_clint_mtime_put = EN_sb_clint_mtime_put ;

  // action method sb_ext_interrupt_put
  assign RDY_sb_ext_interrupt_put = 1'd1 ;
  assign CAN_FIRE_sb_ext_interrupt_put = 1'd1 ;
  assign WILL_FIRE_sb_ext_interrupt_put = EN_sb_ext_interrupt_put ;

  // actionvalue method io_dump_get
  assign io_dump_get =
	     { (riscv_dump_get[166:165] == 2'd3) ?
		 riscv_dump_get[166:165] :
		 2'd0,
	       riscv_dump_get[164:0] } ;
  assign RDY_io_dump_get = riscv_RDY_dump_get ;
  assign CAN_FIRE_io_dump_get = riscv_RDY_dump_get ;
  assign WILL_FIRE_io_dump_get = EN_io_dump_get ;

  // submodule fetch_xactor_f_rd_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) fetch_xactor_f_rd_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(fetch_xactor_f_rd_addr_D_IN),
								  .ENQ(fetch_xactor_f_rd_addr_ENQ),
								  .DEQ(fetch_xactor_f_rd_addr_DEQ),
								  .CLR(fetch_xactor_f_rd_addr_CLR),
								  .D_OUT(fetch_xactor_f_rd_addr_D_OUT),
								  .FULL_N(fetch_xactor_f_rd_addr_FULL_N),
								  .EMPTY_N(fetch_xactor_f_rd_addr_EMPTY_N));

  // submodule fetch_xactor_f_rd_data
  FIFO2 #(.width(32'd66), .guarded(32'd1)) fetch_xactor_f_rd_data(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(fetch_xactor_f_rd_data_D_IN),
								  .ENQ(fetch_xactor_f_rd_data_ENQ),
								  .DEQ(fetch_xactor_f_rd_data_DEQ),
								  .CLR(fetch_xactor_f_rd_data_CLR),
								  .D_OUT(fetch_xactor_f_rd_data_D_OUT),
								  .FULL_N(fetch_xactor_f_rd_data_FULL_N),
								  .EMPTY_N(fetch_xactor_f_rd_data_EMPTY_N));

  // submodule fetch_xactor_f_wr_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) fetch_xactor_f_wr_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(fetch_xactor_f_wr_addr_D_IN),
								  .ENQ(fetch_xactor_f_wr_addr_ENQ),
								  .DEQ(fetch_xactor_f_wr_addr_DEQ),
								  .CLR(fetch_xactor_f_wr_addr_CLR),
								  .D_OUT(fetch_xactor_f_wr_addr_D_OUT),
								  .FULL_N(),
								  .EMPTY_N(fetch_xactor_f_wr_addr_EMPTY_N));

  // submodule fetch_xactor_f_wr_data
  FIFO2 #(.width(32'd72), .guarded(32'd1)) fetch_xactor_f_wr_data(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(fetch_xactor_f_wr_data_D_IN),
								  .ENQ(fetch_xactor_f_wr_data_ENQ),
								  .DEQ(fetch_xactor_f_wr_data_DEQ),
								  .CLR(fetch_xactor_f_wr_data_CLR),
								  .D_OUT(fetch_xactor_f_wr_data_D_OUT),
								  .FULL_N(),
								  .EMPTY_N(fetch_xactor_f_wr_data_EMPTY_N));

  // submodule fetch_xactor_f_wr_resp
  FIFO2 #(.width(32'd2), .guarded(32'd1)) fetch_xactor_f_wr_resp(.RST(RST_N),
								 .CLK(CLK),
								 .D_IN(fetch_xactor_f_wr_resp_D_IN),
								 .ENQ(fetch_xactor_f_wr_resp_ENQ),
								 .DEQ(fetch_xactor_f_wr_resp_DEQ),
								 .CLR(fetch_xactor_f_wr_resp_CLR),
								 .D_OUT(),
								 .FULL_N(fetch_xactor_f_wr_resp_FULL_N),
								 .EMPTY_N());

  // submodule ff_atomic_state
  FIFO1 #(.width(32'd64), .guarded(32'd1)) ff_atomic_state(.RST(RST_N),
							   .CLK(CLK),
							   .D_IN(ff_atomic_state_D_IN),
							   .ENQ(ff_atomic_state_ENQ),
							   .DEQ(ff_atomic_state_DEQ),
							   .CLR(ff_atomic_state_CLR),
							   .D_OUT(ff_atomic_state_D_OUT),
							   .FULL_N(ff_atomic_state_FULL_N),
							   .EMPTY_N(ff_atomic_state_EMPTY_N));

  // submodule ff_inst_access_fault
  FIFO2 #(.width(32'd1), .guarded(32'd1)) ff_inst_access_fault(.RST(RST_N),
							       .CLK(CLK),
							       .D_IN(ff_inst_access_fault_D_IN),
							       .ENQ(ff_inst_access_fault_ENQ),
							       .DEQ(ff_inst_access_fault_DEQ),
							       .CLR(ff_inst_access_fault_CLR),
							       .D_OUT(ff_inst_access_fault_D_OUT),
							       .FULL_N(ff_inst_access_fault_FULL_N),
							       .EMPTY_N(ff_inst_access_fault_EMPTY_N));

  // submodule ff_inst_request
  FIFO2 #(.width(32'd66), .guarded(32'd1)) ff_inst_request(.RST(RST_N),
							   .CLK(CLK),
							   .D_IN(ff_inst_request_D_IN),
							   .ENQ(ff_inst_request_ENQ),
							   .DEQ(ff_inst_request_DEQ),
							   .CLR(ff_inst_request_CLR),
							   .D_OUT(ff_inst_request_D_OUT),
							   .FULL_N(ff_inst_request_FULL_N),
							   .EMPTY_N(ff_inst_request_EMPTY_N));

  // submodule ff_mem_access_fault
  FIFO2 #(.width(32'd1), .guarded(32'd1)) ff_mem_access_fault(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(ff_mem_access_fault_D_IN),
							      .ENQ(ff_mem_access_fault_ENQ),
							      .DEQ(ff_mem_access_fault_DEQ),
							      .CLR(ff_mem_access_fault_CLR),
							      .D_OUT(),
							      .FULL_N(),
							      .EMPTY_N());

  // submodule ff_mem_request
  FIFO2 #(.width(32'd139), .guarded(32'd1)) ff_mem_request(.RST(RST_N),
							   .CLK(CLK),
							   .D_IN(ff_mem_request_D_IN),
							   .ENQ(ff_mem_request_ENQ),
							   .DEQ(ff_mem_request_DEQ),
							   .CLR(ff_mem_request_CLR),
							   .D_OUT(ff_mem_request_D_OUT),
							   .FULL_N(ff_mem_request_FULL_N),
							   .EMPTY_N(ff_mem_request_EMPTY_N));

  // submodule memory_xactor_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) memory_xactor_f_rd_addr(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(memory_xactor_f_rd_addr_D_IN),
						   .ENQ(memory_xactor_f_rd_addr_ENQ),
						   .DEQ(memory_xactor_f_rd_addr_DEQ),
						   .CLR(memory_xactor_f_rd_addr_CLR),
						   .D_OUT(memory_xactor_f_rd_addr_D_OUT),
						   .FULL_N(memory_xactor_f_rd_addr_FULL_N),
						   .EMPTY_N(memory_xactor_f_rd_addr_EMPTY_N));

  // submodule memory_xactor_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) memory_xactor_f_rd_data(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(memory_xactor_f_rd_data_D_IN),
						   .ENQ(memory_xactor_f_rd_data_ENQ),
						   .DEQ(memory_xactor_f_rd_data_DEQ),
						   .CLR(memory_xactor_f_rd_data_CLR),
						   .D_OUT(memory_xactor_f_rd_data_D_OUT),
						   .FULL_N(memory_xactor_f_rd_data_FULL_N),
						   .EMPTY_N(memory_xactor_f_rd_data_EMPTY_N));

  // submodule memory_xactor_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) memory_xactor_f_wr_addr(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(memory_xactor_f_wr_addr_D_IN),
						   .ENQ(memory_xactor_f_wr_addr_ENQ),
						   .DEQ(memory_xactor_f_wr_addr_DEQ),
						   .CLR(memory_xactor_f_wr_addr_CLR),
						   .D_OUT(memory_xactor_f_wr_addr_D_OUT),
						   .FULL_N(memory_xactor_f_wr_addr_FULL_N),
						   .EMPTY_N(memory_xactor_f_wr_addr_EMPTY_N));

  // submodule memory_xactor_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) memory_xactor_f_wr_data(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(memory_xactor_f_wr_data_D_IN),
						   .ENQ(memory_xactor_f_wr_data_ENQ),
						   .DEQ(memory_xactor_f_wr_data_DEQ),
						   .CLR(memory_xactor_f_wr_data_CLR),
						   .D_OUT(memory_xactor_f_wr_data_D_OUT),
						   .FULL_N(memory_xactor_f_wr_data_FULL_N),
						   .EMPTY_N(memory_xactor_f_wr_data_EMPTY_N));

  // submodule memory_xactor_f_wr_resp
  FIFO2 #(.width(32'd2), .guarded(32'd1)) memory_xactor_f_wr_resp(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(memory_xactor_f_wr_resp_D_IN),
								  .ENQ(memory_xactor_f_wr_resp_ENQ),
								  .DEQ(memory_xactor_f_wr_resp_DEQ),
								  .CLR(memory_xactor_f_wr_resp_CLR),
								  .D_OUT(memory_xactor_f_wr_resp_D_OUT),
								  .FULL_N(memory_xactor_f_wr_resp_FULL_N),
								  .EMPTY_N(memory_xactor_f_wr_resp_EMPTY_N));

  // submodule riscv
  mkriscv riscv(.resetpc(resetpc),
		.CLK(CLK),
		.RST_N(RST_N),
		.clint_msip_intrpt(riscv_clint_msip_intrpt),
		.clint_mtime_c_mtime(riscv_clint_mtime_c_mtime),
		.clint_mtip_intrpt(riscv_clint_mtip_intrpt),
		.ext_interrupt_intrpt(riscv_ext_interrupt_intrpt),
		.inst_response_put(riscv_inst_response_put),
		.memory_response_put(riscv_memory_response_put),
		.EN_inst_request_get(riscv_EN_inst_request_get),
		.EN_inst_response_put(riscv_EN_inst_response_put),
		.EN_memory_request_get(riscv_EN_memory_request_get),
		.EN_memory_response_put(riscv_EN_memory_response_put),
		.EN_clint_msip(riscv_EN_clint_msip),
		.EN_clint_mtip(riscv_EN_clint_mtip),
		.EN_clint_mtime(riscv_EN_clint_mtime),
		.EN_ext_interrupt(riscv_EN_ext_interrupt),
		.EN_dump_get(riscv_EN_dump_get),
		.inst_request_get(riscv_inst_request_get),
		.RDY_inst_request_get(riscv_RDY_inst_request_get),
		.RDY_inst_response_put(riscv_RDY_inst_response_put),
		.memory_request_get(riscv_memory_request_get),
		.RDY_memory_request_get(riscv_RDY_memory_request_get),
		.RDY_memory_response_put(),
		.RDY_clint_msip(),
		.RDY_clint_mtip(),
		.RDY_clint_mtime(),
		.RDY_ext_interrupt(),
		.dump_get(riscv_dump_get),
		.RDY_dump_get(riscv_RDY_dump_get),
		.mv_curr_priv(riscv_mv_curr_priv),
		.RDY_mv_curr_priv(),
		.mv_trap(riscv_mv_trap),
		.RDY_mv_trap(),
		.mv_pmp_cfg(riscv_mv_pmp_cfg),
		.RDY_mv_pmp_cfg(),
		.mv_pmp_addr(riscv_mv_pmp_addr),
		.RDY_mv_pmp_addr());

  // rule RL_handle_fetch_request
  assign CAN_FIRE_RL_handle_fetch_request =
	     riscv_RDY_inst_request_get && ff_inst_access_fault_FULL_N &&
	     ff_inst_request_FULL_N &&
	     fetch_xactor_f_rd_addr_FULL_N ;
  assign WILL_FIRE_RL_handle_fetch_request =
	     CAN_FIRE_RL_handle_fetch_request ;

  // rule RL_handle_fetch_response
  assign CAN_FIRE_RL_handle_fetch_response =
	     riscv_RDY_inst_response_put && ff_inst_access_fault_EMPTY_N &&
	     fetch_xactor_f_rd_data_EMPTY_N &&
	     ff_inst_request_EMPTY_N &&
	     !ff_inst_access_fault_D_OUT ;
  assign WILL_FIRE_RL_handle_fetch_response =
	     CAN_FIRE_RL_handle_fetch_response ;

  // rule RL_handle_inst_access_fault
  assign CAN_FIRE_RL_handle_inst_access_fault =
	     riscv_RDY_inst_response_put && ff_inst_access_fault_EMPTY_N &&
	     ff_inst_request_EMPTY_N &&
	     ff_inst_access_fault_D_OUT ;
  assign WILL_FIRE_RL_handle_inst_access_fault =
	     CAN_FIRE_RL_handle_inst_access_fault ;

  // rule RL_handle_memory_request
  assign CAN_FIRE_RL_handle_memory_request =
	     riscv_RDY_memory_request_get && ff_mem_request_FULL_N &&
	     memory_xactor_f_rd_addr_FULL_N &&
	     memory_xactor_f_wr_addr_FULL_N &&
	     memory_xactor_f_wr_data_FULL_N ;
  assign WILL_FIRE_RL_handle_memory_request =
	     CAN_FIRE_RL_handle_memory_request && !riscv_mv_trap ;

  // rule RL_handle_memoryRead_response
  assign CAN_FIRE_RL_handle_memoryRead_response =
	     ff_mem_request_EMPTY_N && memory_xactor_f_rd_data_EMPTY_N &&
	     ff_mem_request_D_OUT[10:9] == 2'd0 ;
  assign WILL_FIRE_RL_handle_memoryRead_response =
	     CAN_FIRE_RL_handle_memoryRead_response ;

  // rule RL_handle_memoryWrite_response
  assign CAN_FIRE_RL_handle_memoryWrite_response =
	     ff_mem_request_EMPTY_N && memory_xactor_f_wr_resp_EMPTY_N &&
	     ff_mem_request_D_OUT[10:9] == 2'd1 ;
  assign WILL_FIRE_RL_handle_memoryWrite_response =
	     CAN_FIRE_RL_handle_memoryWrite_response ;

  // rule RL_handle_atomic_readresponse
  assign CAN_FIRE_RL_handle_atomic_readresponse =
	     ff_mem_request_EMPTY_N && memory_xactor_f_rd_data_EMPTY_N &&
	     memory_xactor_f_wr_addr_FULL_N &&
	     memory_xactor_f_wr_data_FULL_N &&
	     ff_atomic_state_FULL_N &&
	     ff_mem_request_D_OUT[10:9] != 2'd0 &&
	     ff_mem_request_D_OUT[10:9] != 2'd1 &&
	     ff_mem_request_D_OUT[10:9] != 2'd3 &&
	     !ff_atomic_state_EMPTY_N ;
  assign WILL_FIRE_RL_handle_atomic_readresponse =
	     CAN_FIRE_RL_handle_atomic_readresponse &&
	     !WILL_FIRE_RL_handle_memory_request ;

  // rule RL_update_epochs
  assign CAN_FIRE_RL_update_epochs = riscv_mv_trap ;
  assign WILL_FIRE_RL_update_epochs = riscv_mv_trap ;

  // rule RL_handle_atomic_writeresponse
  assign CAN_FIRE_RL_handle_atomic_writeresponse =
	     ff_mem_request_EMPTY_N && memory_xactor_f_wr_resp_EMPTY_N &&
	     ff_atomic_state_EMPTY_N &&
	     ff_mem_request_D_OUT[10:9] != 2'd0 &&
	     ff_mem_request_D_OUT[10:9] != 2'd1 &&
	     ff_mem_request_D_OUT[10:9] != 2'd3 ;
  assign WILL_FIRE_RL_handle_atomic_writeresponse =
	     CAN_FIRE_RL_handle_atomic_writeresponse ;

  // inputs to muxes for submodule ports
  assign MUX_memory_xactor_f_wr_addr_enq_1__SEL_1 =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0 ;
  assign MUX_riscv_memory_response_put_1__SEL_1 =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0 ;
  assign MUX_memory_xactor_f_wr_addr_enq_1__VAL_1 =
	     { ff_mem_request_D_OUT[106:75],
	       aw_awprot__h9129,
	       ff_mem_request_D_OUT[7:6] } ;
  assign MUX_memory_xactor_f_wr_addr_enq_1__VAL_2 =
	     { x__h5078[31:0], 3'd1, riscv_memory_request_get[7:6] } ;
  assign MUX_memory_xactor_f_wr_data_enq_1__VAL_1 =
	     (ff_mem_request_D_OUT[8:6] == 3'd3) ?
	       { wdata__h9103, write_strobe__h8725 } :
	       { wdata___1__h9203, write_strobe___1__h9202 } ;
  assign MUX_memory_xactor_f_wr_data_enq_1__VAL_2 =
	     { w_wdata__h5384, w_wstrb__h5385 } ;
  assign MUX_riscv_inst_response_put_1__VAL_1 =
	     { x__h3633[31:0],
	       ff_inst_request_D_OUT[1:0],
	       fetch_xactor_f_rd_data_D_OUT[65:64] != 2'd0 } ;
  assign MUX_riscv_inst_response_put_1__VAL_2 =
	     { ff_inst_request_D_OUT[33:0], 1'd1 } ;
  assign MUX_riscv_memory_response_put_1__VAL_1 =
	     { ff_mem_request_D_OUT[138:75],
	       memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0,
	       ff_mem_request_D_OUT[5] } ;
  assign MUX_riscv_memory_response_put_1__VAL_2 =
	     { put_data__h7891,
	       memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0,
	       ff_mem_request_D_OUT[5] } ;
  assign MUX_riscv_memory_response_put_1__VAL_3 =
	     { put_data__h8506,
	       memory_xactor_f_wr_resp_D_OUT != 2'd0,
	       ff_mem_request_D_OUT[5] } ;
  assign MUX_riscv_memory_response_put_1__VAL_4 =
	     { put_data__h9976,
	       memory_xactor_f_wr_resp_D_OUT != 2'd0,
	       ff_mem_request_D_OUT[5] } ;

  // register rg_wEpoch
  assign rg_wEpoch_D_IN = x_port1__read__h4086 ;
  assign rg_wEpoch_EN = 1'b1 ;

  // submodule fetch_xactor_f_rd_addr
  assign fetch_xactor_f_rd_addr_D_IN =
	     { riscv_inst_request_get[33:2], aw_awprot__h9129, 2'd2 } ;
  assign fetch_xactor_f_rd_addr_ENQ =
	     WILL_FIRE_RL_handle_fetch_request &&
	     riscv_inst_request_get[65:34] == 32'd0 &&
	     !fn_pmp_lookup___d21[6] ;
  assign fetch_xactor_f_rd_addr_DEQ =
	     fetch_xactor_f_rd_addr_EMPTY_N && master_i_m_arready_arready ;
  assign fetch_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule fetch_xactor_f_rd_data
  assign fetch_xactor_f_rd_data_D_IN =
	     { master_i_m_rvalid_rresp, master_i_m_rvalid_rdata } ;
  assign fetch_xactor_f_rd_data_ENQ =
	     master_i_m_rvalid_rvalid && fetch_xactor_f_rd_data_FULL_N ;
  assign fetch_xactor_f_rd_data_DEQ = CAN_FIRE_RL_handle_fetch_response ;
  assign fetch_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule fetch_xactor_f_wr_addr
  assign fetch_xactor_f_wr_addr_D_IN = 37'h0 ;
  assign fetch_xactor_f_wr_addr_ENQ = 1'b0 ;
  assign fetch_xactor_f_wr_addr_DEQ =
	     fetch_xactor_f_wr_addr_EMPTY_N && master_i_m_awready_awready ;
  assign fetch_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule fetch_xactor_f_wr_data
  assign fetch_xactor_f_wr_data_D_IN = 72'h0 ;
  assign fetch_xactor_f_wr_data_ENQ = 1'b0 ;
  assign fetch_xactor_f_wr_data_DEQ =
	     fetch_xactor_f_wr_data_EMPTY_N && master_i_m_wready_wready ;
  assign fetch_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule fetch_xactor_f_wr_resp
  assign fetch_xactor_f_wr_resp_D_IN = master_i_m_bvalid_bresp ;
  assign fetch_xactor_f_wr_resp_ENQ =
	     master_i_m_bvalid_bvalid && fetch_xactor_f_wr_resp_FULL_N ;
  assign fetch_xactor_f_wr_resp_DEQ = 1'b0 ;
  assign fetch_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule ff_atomic_state
  assign ff_atomic_state_D_IN =
	     IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d218 ;
  assign ff_atomic_state_ENQ = MUX_memory_xactor_f_wr_addr_enq_1__SEL_1 ;
  assign ff_atomic_state_DEQ = CAN_FIRE_RL_handle_atomic_writeresponse ;
  assign ff_atomic_state_CLR = 1'b0 ;

  // submodule ff_inst_access_fault
  assign ff_inst_access_fault_D_IN =
	     riscv_inst_request_get[65:34] != 32'd0 ||
	     fn_pmp_lookup___d21[6] ;
  assign ff_inst_access_fault_ENQ = CAN_FIRE_RL_handle_fetch_request ;
  assign ff_inst_access_fault_DEQ =
	     WILL_FIRE_RL_handle_inst_access_fault ||
	     WILL_FIRE_RL_handle_fetch_response ;
  assign ff_inst_access_fault_CLR = 1'b0 ;

  // submodule ff_inst_request
  assign ff_inst_request_D_IN = riscv_inst_request_get ;
  assign ff_inst_request_ENQ = CAN_FIRE_RL_handle_fetch_request ;
  assign ff_inst_request_DEQ =
	     WILL_FIRE_RL_handle_inst_access_fault ||
	     WILL_FIRE_RL_handle_fetch_response ;
  assign ff_inst_request_CLR = 1'b0 ;

  // submodule ff_mem_access_fault
  assign ff_mem_access_fault_D_IN = 1'b0 ;
  assign ff_mem_access_fault_ENQ = 1'b0 ;
  assign ff_mem_access_fault_DEQ = 1'b0 ;
  assign ff_mem_access_fault_CLR = 1'b0 ;

  // submodule ff_mem_request
  assign ff_mem_request_D_IN =
	     { x__h5078,
	       w_wdata__h5384,
	       CASE_riscvmemory_request_get_BITS_10_TO_9_0_r_ETC__q6,
	       riscv_memory_request_get[8:0] } ;
  assign ff_mem_request_ENQ =
	     WILL_FIRE_RL_handle_memory_request &&
	     rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 ;
  assign ff_mem_request_DEQ =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0 ||
	     WILL_FIRE_RL_handle_atomic_writeresponse ||
	     WILL_FIRE_RL_handle_memoryWrite_response ||
	     WILL_FIRE_RL_handle_memoryRead_response ;
  assign ff_mem_request_CLR = 1'b0 ;

  // submodule memory_xactor_f_rd_addr
  assign memory_xactor_f_rd_addr_D_IN =
	     MUX_memory_xactor_f_wr_addr_enq_1__VAL_2 ;
  assign memory_xactor_f_rd_addr_ENQ =
	     WILL_FIRE_RL_handle_memory_request &&
	     rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	     riscv_memory_request_get[10:9] != 2'd1 ;
  assign memory_xactor_f_rd_addr_DEQ =
	     memory_xactor_f_rd_addr_EMPTY_N && master_d_m_arready_arready ;
  assign memory_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule memory_xactor_f_rd_data
  assign memory_xactor_f_rd_data_D_IN =
	     { master_d_m_rvalid_rresp, master_d_m_rvalid_rdata } ;
  assign memory_xactor_f_rd_data_ENQ =
	     master_d_m_rvalid_rvalid && memory_xactor_f_rd_data_FULL_N ;
  assign memory_xactor_f_rd_data_DEQ =
	     WILL_FIRE_RL_handle_atomic_readresponse ||
	     WILL_FIRE_RL_handle_memoryRead_response ;
  assign memory_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule memory_xactor_f_wr_addr
  assign memory_xactor_f_wr_addr_D_IN =
	     MUX_memory_xactor_f_wr_addr_enq_1__SEL_1 ?
	       MUX_memory_xactor_f_wr_addr_enq_1__VAL_1 :
	       MUX_memory_xactor_f_wr_addr_enq_1__VAL_2 ;
  assign memory_xactor_f_wr_addr_ENQ =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0 ||
	     WILL_FIRE_RL_handle_memory_request &&
	     rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	     riscv_memory_request_get[10:9] == 2'd1 ;
  assign memory_xactor_f_wr_addr_DEQ =
	     memory_xactor_f_wr_addr_EMPTY_N && master_d_m_awready_awready ;
  assign memory_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule memory_xactor_f_wr_data
  assign memory_xactor_f_wr_data_D_IN =
	     MUX_memory_xactor_f_wr_addr_enq_1__SEL_1 ?
	       MUX_memory_xactor_f_wr_data_enq_1__VAL_1 :
	       MUX_memory_xactor_f_wr_data_enq_1__VAL_2 ;
  assign memory_xactor_f_wr_data_ENQ =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0 ||
	     WILL_FIRE_RL_handle_memory_request &&
	     rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	     riscv_memory_request_get[10:9] == 2'd1 ;
  assign memory_xactor_f_wr_data_DEQ =
	     memory_xactor_f_wr_data_EMPTY_N && master_d_m_wready_wready ;
  assign memory_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule memory_xactor_f_wr_resp
  assign memory_xactor_f_wr_resp_D_IN = master_d_m_bvalid_bresp ;
  assign memory_xactor_f_wr_resp_ENQ =
	     master_d_m_bvalid_bvalid && memory_xactor_f_wr_resp_FULL_N ;
  assign memory_xactor_f_wr_resp_DEQ =
	     WILL_FIRE_RL_handle_atomic_writeresponse ||
	     WILL_FIRE_RL_handle_memoryWrite_response ;
  assign memory_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule riscv
  assign riscv_clint_msip_intrpt = sb_clint_msip_put ;
  assign riscv_clint_mtime_c_mtime = sb_clint_mtime_put ;
  assign riscv_clint_mtip_intrpt = sb_clint_mtip_put ;
  assign riscv_ext_interrupt_intrpt = sb_ext_interrupt_put ;
  assign riscv_inst_response_put =
	     WILL_FIRE_RL_handle_fetch_response ?
	       MUX_riscv_inst_response_put_1__VAL_1 :
	       MUX_riscv_inst_response_put_1__VAL_2 ;
  always@(MUX_riscv_memory_response_put_1__SEL_1 or
	  MUX_riscv_memory_response_put_1__VAL_1 or
	  WILL_FIRE_RL_handle_memoryRead_response or
	  MUX_riscv_memory_response_put_1__VAL_2 or
	  WILL_FIRE_RL_handle_memoryWrite_response or
	  MUX_riscv_memory_response_put_1__VAL_3 or
	  WILL_FIRE_RL_handle_atomic_writeresponse or
	  MUX_riscv_memory_response_put_1__VAL_4)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_riscv_memory_response_put_1__SEL_1:
	  riscv_memory_response_put = MUX_riscv_memory_response_put_1__VAL_1;
      WILL_FIRE_RL_handle_memoryRead_response:
	  riscv_memory_response_put = MUX_riscv_memory_response_put_1__VAL_2;
      WILL_FIRE_RL_handle_memoryWrite_response:
	  riscv_memory_response_put = MUX_riscv_memory_response_put_1__VAL_3;
      WILL_FIRE_RL_handle_atomic_writeresponse:
	  riscv_memory_response_put = MUX_riscv_memory_response_put_1__VAL_4;
      default: riscv_memory_response_put =
		   66'h2AAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign riscv_EN_inst_request_get = CAN_FIRE_RL_handle_fetch_request ;
  assign riscv_EN_inst_response_put =
	     WILL_FIRE_RL_handle_fetch_response ||
	     WILL_FIRE_RL_handle_inst_access_fault ;
  assign riscv_EN_memory_request_get = WILL_FIRE_RL_handle_memory_request ;
  assign riscv_EN_memory_response_put =
	     WILL_FIRE_RL_handle_atomic_readresponse &&
	     memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0 ||
	     WILL_FIRE_RL_handle_memoryRead_response ||
	     WILL_FIRE_RL_handle_memoryWrite_response ||
	     WILL_FIRE_RL_handle_atomic_writeresponse ;
  assign riscv_EN_clint_msip = EN_sb_clint_msip_put ;
  assign riscv_EN_clint_mtip = EN_sb_clint_mtip_put ;
  assign riscv_EN_clint_mtime = EN_sb_clint_mtime_put ;
  assign riscv_EN_ext_interrupt = EN_sb_ext_interrupt_put ;
  assign riscv_EN_dump_get = EN_io_dump_get ;

  // remaining internal signals
  module_fn_pmp_lookup instance_fn_pmp_lookup_1(.fn_pmp_lookup_req({ pmpreq_address__h1928,
								     8'd18 }),
						.fn_pmp_lookup_priv(IF_riscv_mv_curr_priv__6_EQ_3_7_THEN_riscv_mv__ETC___d18),
						.fn_pmp_lookup_pmpcfg(riscv_mv_pmp_cfg),
						.fn_pmp_lookup_pmpaddr(riscv_mv_pmp_addr),
						.fn_pmp_lookup(fn_pmp_lookup___d21));
  module_fn_pmp_lookup instance_fn_pmp_lookup_0(.fn_pmp_lookup_req({ pmpreq_address__h4100,
								     pmpreq_num_bytes__h4101,
								     pmpreq_access_type__h4102 }),
						.fn_pmp_lookup_priv(IF_riscv_mv_curr_priv__6_EQ_3_7_THEN_riscv_mv__ETC___d18),
						.fn_pmp_lookup_pmpcfg(riscv_mv_pmp_cfg),
						.fn_pmp_lookup_pmpaddr(riscv_mv_pmp_addr),
						.fn_pmp_lookup(fn_pmp_lookup___d119));
  assign IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d218 =
	     (ff_mem_request_D_OUT[7:6] == 2'd2) ?
	       IF_ff_mem_request_first__90_BIT_8_99_THEN_0_CO_ETC___d217 :
	       rdata__h7865 ;
  assign IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC__q3 =
	     IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d218[31:0] ;
  assign IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d317 =
	     op1__h9481 <= op2__h9482 ;
  assign IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d322 =
	     (op1__h9481 ^ 64'h8000000000000000) <=
	     (op2__h9482 ^ 64'h8000000000000000) ;
  assign IF_ff_mem_request_first__90_BIT_8_99_THEN_0_CO_ETC___d217 =
	     ff_mem_request_D_OUT[8] ?
	       { 32'd0, rdata__h7865[31:0] } :
	       { {32{rdata865_BITS_31_TO_0__q2[31]}},
		 rdata865_BITS_31_TO_0__q2 } ;
  assign IF_riscv_mv_curr_priv__6_EQ_3_7_THEN_riscv_mv__ETC___d18 =
	     (riscv_mv_curr_priv == 2'd3) ? riscv_mv_curr_priv : 2'd0 ;
  assign aw_awprot__h9129 = { 2'd0, riscv_mv_curr_priv[1] } ;
  assign ff_mem_requestD_OUT_BITS_42_TO_11__q1 = ff_mem_request_D_OUT[42:11] ;
  assign lv_data__h3600 =
	     fetch_xactor_f_rd_data_D_OUT[63:0] >> lv_shift__h3599 ;
  assign lv_shift__h3599 = { ff_inst_request_D_OUT[4:2], 3'd0 } ;
  assign lv_shift__h7864 = { ff_mem_request_D_OUT[77:75], 3'd0 } ;
  assign op1___1__h9539 =
	     { {32{IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC__q3[31]}},
	       IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC__q3 } ;
  assign op1__h9481 =
	     ff_mem_request_D_OUT[4] ?
	       IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d218 :
	       op1___1__h9539 ;
  assign op2___1__h9540 =
	     { {32{ff_mem_requestD_OUT_BITS_42_TO_11__q1[31]}},
	       ff_mem_requestD_OUT_BITS_42_TO_11__q1 } ;
  assign op2__h9482 =
	     ff_mem_request_D_OUT[4] ?
	       ff_mem_request_D_OUT[74:11] :
	       op2___1__h9540 ;
  assign pmpreq_access_type__h4102 =
	     (riscv_memory_request_get[10:9] == 2'd0) ?
	       riscv_memory_request_get[10:9] :
	       2'd1 ;
  assign pmpreq_address__h1928 = riscv_inst_request_get[33:2] ;
  assign pmpreq_address__h4100 = riscv_memory_request_get[106:75] ;
  assign pmpreq_num_bytes__h4101 = { 4'd0, riscv_memory_request_get[7:6] } ;
  assign put_data__h7891 =
	     (memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0) ?
	       IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220 :
	       ff_mem_request_D_OUT[138:75] ;
  assign put_data__h8506 =
	     (memory_xactor_f_wr_resp_D_OUT == 2'd0) ?
	       64'd0 :
	       ff_mem_request_D_OUT[138:75] ;
  assign put_data__h9976 =
	     (memory_xactor_f_wr_resp_D_OUT == 2'd0) ?
	       ff_atomic_state_D_OUT :
	       ff_mem_request_D_OUT[138:75] ;
  assign rdata865_BITS_15_TO_0__q5 = rdata__h7865[15:0] ;
  assign rdata865_BITS_31_TO_0__q2 = rdata__h7865[31:0] ;
  assign rdata865_BITS_7_TO_0__q4 = rdata__h7865[7:0] ;
  assign rdata__h7865 =
	     memory_xactor_f_rd_data_D_OUT[63:0] >> lv_shift__h7864 ;
  assign rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 =
	     x_port1__read__h4086 == riscv_memory_request_get[5] ;
  assign w_wstrb__h5385 =
	     (riscv_memory_request_get[8:6] == 3'd3) ?
	       write_strobe__h4071 :
	       write_strobe___1__h7282 ;
  assign wdata___1__h9203 = {2{wdata__h9103[31:0]}} ;
  assign write_strobe___1__h7282 =
	     write_strobe__h4071 << riscv_memory_request_get[77:75] ;
  assign write_strobe___1__h9202 =
	     write_strobe__h8725 << ff_mem_request_D_OUT[77:75] ;
  assign write_strobe__h8725 =
	     (ff_mem_request_D_OUT[8:6] == 3'd2) ? 8'h0F : 8'd255 ;
  assign x__h3633 =
	     (fetch_xactor_f_rd_data_D_OUT[65:64] == 2'd0) ?
	       lv_data__h3600 :
	       ff_inst_request_D_OUT[65:2] ;
  assign x__h5078 =
	     fn_pmp_lookup___d119[6] ?
	       64'd0 :
	       riscv_memory_request_get[138:75] ;
  assign x_port1__read__h4086 = riscv_mv_trap ? ~rg_wEpoch : rg_wEpoch ;
  always@(riscv_memory_request_get)
  begin
    case (riscv_memory_request_get[7:6])
      2'd0: w_wdata__h5384 = {8{riscv_memory_request_get[18:11]}};
      2'd1: w_wdata__h5384 = {4{riscv_memory_request_get[26:11]}};
      2'd2: w_wdata__h5384 = {2{riscv_memory_request_get[42:11]}};
      2'd3: w_wdata__h5384 = riscv_memory_request_get[74:11];
    endcase
  end
  always@(riscv_memory_request_get)
  begin
    case (riscv_memory_request_get[8:6])
      3'd0: write_strobe__h4071 = 8'b00000001;
      3'd1: write_strobe__h4071 = 8'b00000011;
      3'd2: write_strobe__h4071 = 8'h0F;
      default: write_strobe__h4071 = 8'd255;
    endcase
  end
  always@(ff_mem_request_D_OUT or
	  rdata__h7865 or
	  rdata865_BITS_7_TO_0__q4 or
	  rdata865_BITS_15_TO_0__q5 or
	  IF_ff_mem_request_first__90_BIT_8_99_THEN_0_CO_ETC___d217)
  begin
    case (ff_mem_request_D_OUT[7:6])
      2'd0:
	  IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220 =
	      ff_mem_request_D_OUT[8] ?
		{ 56'd0, rdata__h7865[7:0] } :
		{ {56{rdata865_BITS_7_TO_0__q4[7]}},
		  rdata865_BITS_7_TO_0__q4 };
      2'd1:
	  IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220 =
	      ff_mem_request_D_OUT[8] ?
		{ 48'd0, rdata__h7865[15:0] } :
		{ {48{rdata865_BITS_15_TO_0__q5[15]}},
		  rdata865_BITS_15_TO_0__q5 };
      2'd2:
	  IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220 =
	      IF_ff_mem_request_first__90_BIT_8_99_THEN_0_CO_ETC___d217;
      2'd3:
	  IF_ff_mem_request_first__90_BITS_7_TO_6_97_EQ__ETC___d220 =
	      rdata__h7865;
    endcase
  end
  always@(ff_mem_request_D_OUT or
	  op1__h9481 or
	  op2__h9482 or
	  IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d322 or
	  IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d317)
  begin
    case (ff_mem_request_D_OUT[3:0])
      4'b0: wdata__h9103 = op1__h9481 + op2__h9482;
      4'b0010: wdata__h9103 = op1__h9481 ^ op2__h9482;
      4'b0011: wdata__h9103 = op2__h9482;
      4'b0100: wdata__h9103 = op1__h9481 | op2__h9482;
      4'b0110: wdata__h9103 = op1__h9481 & op2__h9482;
      4'b1000:
	  wdata__h9103 =
	      IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d322 ?
		op1__h9481 :
		op2__h9482;
      4'b1010:
	  wdata__h9103 =
	      IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d322 ?
		op2__h9482 :
		op1__h9481;
      4'b1100:
	  wdata__h9103 =
	      IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d317 ?
		op1__h9481 :
		op2__h9482;
      4'b1110:
	  wdata__h9103 =
	      IF_ff_mem_request_first__90_BIT_4_00_THEN_IF_f_ETC___d317 ?
		op2__h9482 :
		op1__h9481;
      default: wdata__h9103 = op1__h9481;
    endcase
  end
  always@(riscv_memory_request_get)
  begin
    case (riscv_memory_request_get[10:9])
      2'd0, 2'd1, 2'd3:
	  CASE_riscvmemory_request_get_BITS_10_TO_9_0_r_ETC__q6 =
	      riscv_memory_request_get[10:9];
      2'd2: CASE_riscvmemory_request_get_BITS_10_TO_9_0_r_ETC__q6 = 2'd2;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_wEpoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_wEpoch_EN) rg_wEpoch <= `BSV_ASSIGNMENT_DELAY rg_wEpoch_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_wEpoch = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get[65:34] == 32'd0 &&
	  !fn_pmp_lookup___d21[6])
	begin
	  TASK_testplusargs___d28 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get[65:34] == 32'd0 &&
	  !fn_pmp_lookup___d21[6])
	begin
	  TASK_testplusargs___d29 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get[65:34] == 32'd0 &&
	  !fn_pmp_lookup___d21[6])
	begin
	  TASK_testplusargs___d30 = $test$plusargs("l0");
	  #0;
	end
    riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33 =
	riscv_inst_request_get[65:34] == 32'd0 && !fn_pmp_lookup___d21[6] &&
	(TASK_testplusargs___d28 ||
	 TASK_testplusargs___d29 && TASK_testplusargs___d30);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get[65:34] == 32'd0 &&
	  !fn_pmp_lookup___d21[6])
	begin
	  v__h3195 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("[%10d", v__h3195, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("CORE : Fetch Request ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("AXI4_Lite_Rd_Addr { ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("'h%h", riscv_inst_request_get[33:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("'h%h", 1'b0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("'h%h", aw_awprot__h9129);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("'h%h", 2'd2, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  riscv_inst_request_get_1_BITS_65_TO_34_2_EQ_0__ETC___d33)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  (riscv_inst_request_get[65:34] != 32'd0 || fn_pmp_lookup___d21[6]))
	begin
	  TASK_testplusargs___d37 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  (riscv_inst_request_get[65:34] != 32'd0 || fn_pmp_lookup___d21[6]))
	begin
	  TASK_testplusargs___d38 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  (riscv_inst_request_get[65:34] != 32'd0 || fn_pmp_lookup___d21[6]))
	begin
	  TASK_testplusargs___d39 = $test$plusargs("l0");
	  #0;
	end
    NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42 =
	(riscv_inst_request_get[65:34] != 32'd0 || fn_pmp_lookup___d21[6]) &&
	(TASK_testplusargs___d37 ||
	 TASK_testplusargs___d38 && TASK_testplusargs___d39);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  (riscv_inst_request_get[65:34] != 32'd0 || fn_pmp_lookup___d21[6]))
	begin
	  v__h3370 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("[%10d", v__h3370, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("CORE : Fetch Request is Faulty: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("InstRequest { ", "addr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("'h%h", riscv_inst_request_get[65:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write(", ", "epoch: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("'h%h", riscv_inst_request_get[1:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_request &&
	  NOT_riscv_inst_request_get_1_BITS_65_TO_34_2_E_ETC___d42)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response)
	begin
	  TASK_testplusargs___d70 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response)
	begin
	  TASK_testplusargs___d71 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response)
	begin
	  TASK_testplusargs___d72 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d76 =
	(TASK_testplusargs___d70 ||
	 TASK_testplusargs___d71 && TASK_testplusargs___d72) &&
	fetch_xactor_f_rd_data_D_OUT[65:64] == 2'd0;
    TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d78 =
	(TASK_testplusargs___d70 ||
	 TASK_testplusargs___d71 && TASK_testplusargs___d72) &&
	fetch_xactor_f_rd_data_D_OUT[65:64] == 2'd1;
    TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d80 =
	(TASK_testplusargs___d70 ||
	 TASK_testplusargs___d71 && TASK_testplusargs___d72) &&
	fetch_xactor_f_rd_data_D_OUT[65:64] == 2'd2;
    TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d85 =
	(TASK_testplusargs___d70 ||
	 TASK_testplusargs___d71 && TASK_testplusargs___d72) &&
	fetch_xactor_f_rd_data_D_OUT[65:64] != 2'd0 &&
	fetch_xactor_f_rd_data_D_OUT[65:64] != 2'd1 &&
	fetch_xactor_f_rd_data_D_OUT[65:64] != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response)
	begin
	  v__h3802 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("[%10d", v__h3802, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("CORE : Fetch Response ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("AXI4_Lite_Rd_Data { ", "rresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d76)
	$write("AXI4_LITE_OKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d78)
	$write("AXI4_LITE_EXOKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d80)
	$write("AXI4_LITE_SLVERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  TASK_testplusargs_0_OR_TASK_testplusargs_1_AND_ETC___d85)
	$write("AXI4_LITE_DECERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write(", ", "rdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("'h%h", fetch_xactor_f_rd_data_D_OUT[63:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write(", ", "ruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_fetch_response &&
	  (TASK_testplusargs___d70 ||
	   TASK_testplusargs___d71 && TASK_testplusargs___d72))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault)
	begin
	  TASK_testplusargs___d91 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault)
	begin
	  TASK_testplusargs___d92 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault)
	begin
	  TASK_testplusargs___d93 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault)
	begin
	  v__h4000 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault &&
	  (TASK_testplusargs___d91 ||
	   TASK_testplusargs___d92 && TASK_testplusargs___d93))
	$write("[%10d", v__h4000, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault &&
	  (TASK_testplusargs___d91 ||
	   TASK_testplusargs___d92 && TASK_testplusargs___d93))
	$write("CORE : Fetch Access Fault ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_inst_access_fault &&
	  (TASK_testplusargs___d91 ||
	   TASK_testplusargs___d92 && TASK_testplusargs___d93))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d154 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d155 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d156 = $test$plusargs("l0 ");
	  #0;
	end
    riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159 =
	riscv_memory_request_get[10:9] == 2'd1 &&
	(TASK_testplusargs___d154 ||
	 TASK_testplusargs___d155 && TASK_testplusargs___d156);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  v__h7409 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("[%10d", v__h7409, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("CORE : Memory write Request ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("AXI4_Lite_Wr_Addr { ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("'h%h", x__h5078[31:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("'h%h", 1'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("'h%h", 3'd1);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("'h%h", riscv_memory_request_get[7:6], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d159)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d162 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d163 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  TASK_testplusargs___d164 = $test$plusargs("l0 ");
	  #0;
	end
    riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167 =
	riscv_memory_request_get[10:9] == 2'd1 &&
	(TASK_testplusargs___d162 ||
	 TASK_testplusargs___d163 && TASK_testplusargs___d164);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] == 2'd1)
	begin
	  v__h7569 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("[%10d", v__h7569, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("CORE : Memory write Request ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("AXI4_Lite_Wr_Data { ", "wdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("'h%h", w_wdata__h5384);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write(", ", "wstrb: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("'h%h", w_wstrb__h5385, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get_07_BITS_10_TO_9_10_EQ_ETC___d167)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] != 2'd1)
	begin
	  TASK_testplusargs___d172 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] != 2'd1)
	begin
	  TASK_testplusargs___d173 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] != 2'd1)
	begin
	  TASK_testplusargs___d174 = $test$plusargs("l0");
	  #0;
	end
    NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177 =
	riscv_memory_request_get[10:9] != 2'd1 &&
	(TASK_testplusargs___d172 ||
	 TASK_testplusargs___d173 && TASK_testplusargs___d174);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  riscv_memory_request_get[10:9] != 2'd1)
	begin
	  v__h5179 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("[%10d", v__h5179, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("CORE : Memory Read Request ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("AXI4_Lite_Rd_Addr { ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("'h%h", x__h5078[31:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("'h%h", 1'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("'h%h", 3'd1);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("'h%h", riscv_memory_request_get[7:6], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memory_request &&
	  rg_wEpoch_port1__read__06_EQ_riscv_memory_requ_ETC___d109 &&
	  NOT_riscv_memory_request_get_07_BITS_10_TO_9_1_ETC___d177)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response)
	begin
	  TASK_testplusargs___d227 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response)
	begin
	  TASK_testplusargs___d228 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response)
	begin
	  TASK_testplusargs___d229 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d233 =
	(TASK_testplusargs___d227 ||
	 TASK_testplusargs___d228 && TASK_testplusargs___d229) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0;
    TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d235 =
	(TASK_testplusargs___d227 ||
	 TASK_testplusargs___d228 && TASK_testplusargs___d229) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd1;
    TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d237 =
	(TASK_testplusargs___d227 ||
	 TASK_testplusargs___d228 && TASK_testplusargs___d229) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd2;
    TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d242 =
	(TASK_testplusargs___d227 ||
	 TASK_testplusargs___d228 && TASK_testplusargs___d229) &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0 &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd1 &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response)
	begin
	  v__h8304 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("[%10d", v__h8304, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("CORE : Memory Read Response ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("AXI4_Lite_Rd_Data { ", "rresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d233)
	$write("AXI4_LITE_OKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d235)
	$write("AXI4_LITE_EXOKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d237)
	$write("AXI4_LITE_SLVERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  TASK_testplusargs_27_OR_TASK_testplusargs_28_A_ETC___d242)
	$write("AXI4_LITE_DECERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write(", ", "rdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("'h%h", memory_xactor_f_rd_data_D_OUT[63:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write(", ", "ruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryRead_response &&
	  (TASK_testplusargs___d227 ||
	   TASK_testplusargs___d228 && TASK_testplusargs___d229))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response)
	begin
	  TASK_testplusargs___d253 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response)
	begin
	  TASK_testplusargs___d254 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response)
	begin
	  TASK_testplusargs___d255 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d259 =
	(TASK_testplusargs___d253 ||
	 TASK_testplusargs___d254 && TASK_testplusargs___d255) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd0;
    TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d261 =
	(TASK_testplusargs___d253 ||
	 TASK_testplusargs___d254 && TASK_testplusargs___d255) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd1;
    TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d263 =
	(TASK_testplusargs___d253 ||
	 TASK_testplusargs___d254 && TASK_testplusargs___d255) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd2;
    TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d268 =
	(TASK_testplusargs___d253 ||
	 TASK_testplusargs___d254 && TASK_testplusargs___d255) &&
	memory_xactor_f_wr_resp_D_OUT != 2'd0 &&
	memory_xactor_f_wr_resp_D_OUT != 2'd1 &&
	memory_xactor_f_wr_resp_D_OUT != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response)
	begin
	  v__h8610 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write("[%10d", v__h8610, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write("CORE : Memory Write Response ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write("AXI4_Lite_Wr_Resp { ", "bresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d259)
	$write("AXI4_LITE_OKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d261)
	$write("AXI4_LITE_EXOKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d263)
	$write("AXI4_LITE_SLVERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  TASK_testplusargs_53_OR_TASK_testplusargs_54_A_ETC___d268)
	$write("AXI4_LITE_DECERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write(", ", "buser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_memoryWrite_response &&
	  (TASK_testplusargs___d253 ||
	   TASK_testplusargs___d254 && TASK_testplusargs___d255))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse)
	begin
	  TASK_testplusargs___d284 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse)
	begin
	  TASK_testplusargs___d285 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse)
	begin
	  TASK_testplusargs___d286 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d290 =
	(TASK_testplusargs___d284 ||
	 TASK_testplusargs___d285 && TASK_testplusargs___d286) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd0;
    TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d291 =
	(TASK_testplusargs___d284 ||
	 TASK_testplusargs___d285 && TASK_testplusargs___d286) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd1;
    TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d292 =
	(TASK_testplusargs___d284 ||
	 TASK_testplusargs___d285 && TASK_testplusargs___d286) &&
	memory_xactor_f_rd_data_D_OUT[65:64] == 2'd2;
    TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d293 =
	(TASK_testplusargs___d284 ||
	 TASK_testplusargs___d285 && TASK_testplusargs___d286) &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd0 &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd1 &&
	memory_xactor_f_rd_data_D_OUT[65:64] != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse)
	begin
	  v__h8793 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("[%10d", v__h8793, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("CORE : Atomic Read Response ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("AXI4_Lite_Rd_Data { ", "rresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d290)
	$write("AXI4_LITE_OKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d291)
	$write("AXI4_LITE_EXOKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d292)
	$write("AXI4_LITE_SLVERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  TASK_testplusargs_84_OR_TASK_testplusargs_85_A_ETC___d293)
	$write("AXI4_LITE_DECERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write(", ", "rdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("'h%h", memory_xactor_f_rd_data_D_OUT[63:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write(", ", "ruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_readresponse &&
	  (TASK_testplusargs___d284 ||
	   TASK_testplusargs___d285 && TASK_testplusargs___d286))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse)
	begin
	  TASK_testplusargs___d351 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse)
	begin
	  TASK_testplusargs___d352 = $test$plusargs("meclass");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse)
	begin
	  TASK_testplusargs___d353 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d357 =
	(TASK_testplusargs___d351 ||
	 TASK_testplusargs___d352 && TASK_testplusargs___d353) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd0;
    TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d358 =
	(TASK_testplusargs___d351 ||
	 TASK_testplusargs___d352 && TASK_testplusargs___d353) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd1;
    TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d359 =
	(TASK_testplusargs___d351 ||
	 TASK_testplusargs___d352 && TASK_testplusargs___d353) &&
	memory_xactor_f_wr_resp_D_OUT == 2'd2;
    TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d360 =
	(TASK_testplusargs___d351 ||
	 TASK_testplusargs___d352 && TASK_testplusargs___d353) &&
	memory_xactor_f_wr_resp_D_OUT != 2'd0 &&
	memory_xactor_f_wr_resp_D_OUT != 2'd1 &&
	memory_xactor_f_wr_resp_D_OUT != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse)
	begin
	  v__h10105 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write("[%10d", v__h10105, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write("CORE : Atomic Write Response ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write("AXI4_Lite_Wr_Resp { ", "bresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d357)
	$write("AXI4_LITE_OKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d358)
	$write("AXI4_LITE_EXOKAY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d359)
	$write("AXI4_LITE_SLVERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  TASK_testplusargs_51_OR_TASK_testplusargs_52_A_ETC___d360)
	$write("AXI4_LITE_DECERR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write(", ", "buser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_handle_atomic_writeresponse &&
	  (TASK_testplusargs___d351 ||
	   TASK_testplusargs___d352 && TASK_testplusargs___d353))
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkeclass_axi4lite

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:55:06 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// rvfi_valid                     O     1 const
// rvfi_order                     O    64 const
// rvfi_insn                      O    32 const
// rvfi_trap                      O     1 const
// rvfi_halt                      O     1 const
// rvfi_intr                      O     1 const
// rvfi_mode                      O     2 const
// rvfi_ixl                       O     2 const
// rvfi_mem_addr                  O    32 const
// rvfi_mem_rmask                 O     4 const
// rvfi_mem_wmask                 O     4 const
// rvfi_mem_rdata                 O    32 const
// rvfi_mem_wdata                 O    32 const
// rvfi_rs1_addr                  O     5 const
// rvfi_rs2_addr                  O     5 const
// rvfi_rs1_rdata                 O    32 const
// rvfi_rs2_rdata                 O    32 const
// rvfi_rd_addr                   O     5 const
// rvfi_rd_wdata                  O    32 const
// rvfi_pc_rdata                  O    32 const
// rvfi_pc_wdata                  O    32 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkFormalWrapper(CLK,
		       RST_N,

		       rvfi_valid,

		       rvfi_order,

		       rvfi_insn,

		       rvfi_trap,

		       rvfi_halt,

		       rvfi_intr,

		       rvfi_mode,

		       rvfi_ixl,

		       rvfi_mem_addr,

		       rvfi_mem_rmask,

		       rvfi_mem_wmask,

		       rvfi_mem_rdata,

		       rvfi_mem_wdata,

		       rvfi_rs1_addr,

		       rvfi_rs2_addr,

		       rvfi_rs1_rdata,

		       rvfi_rs2_rdata,

		       rvfi_rd_addr,

		       rvfi_rd_wdata,

		       rvfi_pc_rdata,

		       rvfi_pc_wdata);
  input  CLK;
  input  RST_N;

  // value method rvfi_valid
  output rvfi_valid;

  // value method rvfi_order
  output [63 : 0] rvfi_order;

  // value method rvfi_insn
  output [31 : 0] rvfi_insn;

  // value method rvfi_trap
  output rvfi_trap;

  // value method rvfi_halt
  output rvfi_halt;

  // value method rvfi_intr
  output rvfi_intr;

  // value method rvfi_mode
  output [1 : 0] rvfi_mode;

  // value method rvfi_ixl
  output [1 : 0] rvfi_ixl;

  // value method rvfi_mem_addr
  output [31 : 0] rvfi_mem_addr;

  // value method rvfi_mem_rmask
  output [3 : 0] rvfi_mem_rmask;

  // value method rvfi_mem_wmask
  output [3 : 0] rvfi_mem_wmask;

  // value method rvfi_mem_rdata
  output [31 : 0] rvfi_mem_rdata;

  // value method rvfi_mem_wdata
  output [31 : 0] rvfi_mem_wdata;

  // value method rvfi_rs1_addr
  output [4 : 0] rvfi_rs1_addr;

  // value method rvfi_rs2_addr
  output [4 : 0] rvfi_rs2_addr;

  // value method rvfi_rs1_rdata
  output [31 : 0] rvfi_rs1_rdata;

  // value method rvfi_rs2_rdata
  output [31 : 0] rvfi_rs2_rdata;

  // value method rvfi_rd_addr
  output [4 : 0] rvfi_rd_addr;

  // value method rvfi_rd_wdata
  output [31 : 0] rvfi_rd_wdata;

  // value method rvfi_pc_rdata
  output [31 : 0] rvfi_pc_rdata;

  // value method rvfi_pc_wdata
  output [31 : 0] rvfi_pc_wdata;

  // signals for module outputs
  wire [63 : 0] rvfi_order;
  wire [31 : 0] rvfi_insn,
		rvfi_mem_addr,
		rvfi_mem_rdata,
		rvfi_mem_wdata,
		rvfi_pc_rdata,
		rvfi_pc_wdata,
		rvfi_rd_wdata,
		rvfi_rs1_rdata,
		rvfi_rs2_rdata;
  wire [4 : 0] rvfi_rd_addr, rvfi_rs1_addr, rvfi_rs2_addr;
  wire [3 : 0] rvfi_mem_rmask, rvfi_mem_wmask;
  wire [1 : 0] rvfi_ixl, rvfi_mode;
  wire rvfi_halt, rvfi_intr, rvfi_trap, rvfi_valid;

  // inlined wires
  wire [3 : 0] soc_uart_user_ifc_wr_status_wget;
  wire soc_clint_clint_wr_mtimecmp_written_whas,
       soc_uart_user_ifc_uart_fifoRecv_r_deq_whas,
       soc_uart_user_ifc_uart_fifoXmit_r_enq_whas,
       soc_uart_user_ifc_uart_pwRecvCellCountReset_whas,
       soc_uart_user_ifc_uart_pwRecvEnableBitCount_whas,
       soc_uart_user_ifc_uart_pwRecvResetBitCount_whas,
       soc_uart_user_ifc_uart_pwXmitCellCountReset_whas,
       soc_uart_user_ifc_uart_pwXmitEnableBitCount_whas,
       soc_uart_user_ifc_uart_pwXmitLoadBuffer_whas;

  // register soc_clint_clint_msip
  reg soc_clint_clint_msip;
  wire soc_clint_clint_msip_D_IN, soc_clint_clint_msip_EN;

  // register soc_clint_clint_mtip
  reg soc_clint_clint_mtip;
  wire soc_clint_clint_mtip_D_IN, soc_clint_clint_mtip_EN;

  // register soc_clint_clint_rg_tick
  reg [3 : 0] soc_clint_clint_rg_tick;
  wire [3 : 0] soc_clint_clint_rg_tick_D_IN;
  wire soc_clint_clint_rg_tick_EN;

  // register soc_clint_clint_rgmtime
  reg [63 : 0] soc_clint_clint_rgmtime;
  wire [63 : 0] soc_clint_clint_rgmtime_D_IN;
  wire soc_clint_clint_rgmtime_EN;

  // register soc_clint_clint_rgmtimecmp
  reg [63 : 0] soc_clint_clint_rgmtimecmp;
  wire [63 : 0] soc_clint_clint_rgmtimecmp_D_IN;
  wire soc_clint_clint_rgmtimecmp_EN;

  // register soc_uart_user_ifc_baud_value
  reg [15 : 0] soc_uart_user_ifc_baud_value;
  wire [15 : 0] soc_uart_user_ifc_baud_value_D_IN;
  wire soc_uart_user_ifc_baud_value_EN;

  // register soc_uart_user_ifc_uart_fifoRecv_countReg
  reg [4 : 0] soc_uart_user_ifc_uart_fifoRecv_countReg;
  wire [4 : 0] soc_uart_user_ifc_uart_fifoRecv_countReg_D_IN;
  wire soc_uart_user_ifc_uart_fifoRecv_countReg_EN;

  // register soc_uart_user_ifc_uart_fifoXmit_countReg
  reg [4 : 0] soc_uart_user_ifc_uart_fifoXmit_countReg;
  wire [4 : 0] soc_uart_user_ifc_uart_fifoXmit_countReg_D_IN;
  wire soc_uart_user_ifc_uart_fifoXmit_countReg_EN;

  // register soc_uart_user_ifc_uart_rRecvBitCount
  reg [3 : 0] soc_uart_user_ifc_uart_rRecvBitCount;
  wire [3 : 0] soc_uart_user_ifc_uart_rRecvBitCount_D_IN;
  wire soc_uart_user_ifc_uart_rRecvBitCount_EN;

  // register soc_uart_user_ifc_uart_rRecvCellCount
  reg [3 : 0] soc_uart_user_ifc_uart_rRecvCellCount;
  wire [3 : 0] soc_uart_user_ifc_uart_rRecvCellCount_D_IN;
  wire soc_uart_user_ifc_uart_rRecvCellCount_EN;

  // register soc_uart_user_ifc_uart_rRecvData
  reg soc_uart_user_ifc_uart_rRecvData;
  wire soc_uart_user_ifc_uart_rRecvData_D_IN,
       soc_uart_user_ifc_uart_rRecvData_EN;

  // register soc_uart_user_ifc_uart_rRecvParity
  reg soc_uart_user_ifc_uart_rRecvParity;
  wire soc_uart_user_ifc_uart_rRecvParity_D_IN,
       soc_uart_user_ifc_uart_rRecvParity_EN;

  // register soc_uart_user_ifc_uart_rRecvState
  reg [2 : 0] soc_uart_user_ifc_uart_rRecvState;
  reg [2 : 0] soc_uart_user_ifc_uart_rRecvState_D_IN;
  wire soc_uart_user_ifc_uart_rRecvState_EN;

  // register soc_uart_user_ifc_uart_rXmitBitCount
  reg [3 : 0] soc_uart_user_ifc_uart_rXmitBitCount;
  wire [3 : 0] soc_uart_user_ifc_uart_rXmitBitCount_D_IN;
  wire soc_uart_user_ifc_uart_rXmitBitCount_EN;

  // register soc_uart_user_ifc_uart_rXmitCellCount
  reg [3 : 0] soc_uart_user_ifc_uart_rXmitCellCount;
  wire [3 : 0] soc_uart_user_ifc_uart_rXmitCellCount_D_IN;
  wire soc_uart_user_ifc_uart_rXmitCellCount_EN;

  // register soc_uart_user_ifc_uart_rXmitDataOut
  reg soc_uart_user_ifc_uart_rXmitDataOut;
  reg soc_uart_user_ifc_uart_rXmitDataOut_D_IN;
  wire soc_uart_user_ifc_uart_rXmitDataOut_EN;

  // register soc_uart_user_ifc_uart_rXmitParity
  reg soc_uart_user_ifc_uart_rXmitParity;
  wire soc_uart_user_ifc_uart_rXmitParity_D_IN,
       soc_uart_user_ifc_uart_rXmitParity_EN;

  // register soc_uart_user_ifc_uart_rXmitState
  reg [2 : 0] soc_uart_user_ifc_uart_rXmitState;
  reg [2 : 0] soc_uart_user_ifc_uart_rXmitState_D_IN;
  wire soc_uart_user_ifc_uart_rXmitState_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_0
  reg soc_uart_user_ifc_uart_vrRecvBuffer_0;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_0_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_0_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_1
  reg soc_uart_user_ifc_uart_vrRecvBuffer_1;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_1_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_1_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_2
  reg soc_uart_user_ifc_uart_vrRecvBuffer_2;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_2_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_2_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_3
  reg soc_uart_user_ifc_uart_vrRecvBuffer_3;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_3_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_3_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_4
  reg soc_uart_user_ifc_uart_vrRecvBuffer_4;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_4_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_4_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_5
  reg soc_uart_user_ifc_uart_vrRecvBuffer_5;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_5_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_5_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_6
  reg soc_uart_user_ifc_uart_vrRecvBuffer_6;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_6_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_6_EN;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_7
  reg soc_uart_user_ifc_uart_vrRecvBuffer_7;
  wire soc_uart_user_ifc_uart_vrRecvBuffer_7_D_IN,
       soc_uart_user_ifc_uart_vrRecvBuffer_7_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_0
  reg soc_uart_user_ifc_uart_vrXmitBuffer_0;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_0_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_0_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_1
  reg soc_uart_user_ifc_uart_vrXmitBuffer_1;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_1_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_1_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_2
  reg soc_uart_user_ifc_uart_vrXmitBuffer_2;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_2_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_2_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_3
  reg soc_uart_user_ifc_uart_vrXmitBuffer_3;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_3_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_3_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_4
  reg soc_uart_user_ifc_uart_vrXmitBuffer_4;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_4_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_4_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_5
  reg soc_uart_user_ifc_uart_vrXmitBuffer_5;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_5_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_5_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_6
  reg soc_uart_user_ifc_uart_vrXmitBuffer_6;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_6_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_6_EN;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_7
  reg soc_uart_user_ifc_uart_vrXmitBuffer_7;
  wire soc_uart_user_ifc_uart_vrXmitBuffer_7_D_IN,
       soc_uart_user_ifc_uart_vrXmitBuffer_7_EN;

  // ports of submodule soc_clint_s_xactor_f_rd_addr
  wire [36 : 0] soc_clint_s_xactor_f_rd_addr_D_IN,
		soc_clint_s_xactor_f_rd_addr_D_OUT;
  wire soc_clint_s_xactor_f_rd_addr_CLR,
       soc_clint_s_xactor_f_rd_addr_DEQ,
       soc_clint_s_xactor_f_rd_addr_EMPTY_N,
       soc_clint_s_xactor_f_rd_addr_ENQ,
       soc_clint_s_xactor_f_rd_addr_FULL_N;

  // ports of submodule soc_clint_s_xactor_f_rd_data
  wire [65 : 0] soc_clint_s_xactor_f_rd_data_D_IN,
		soc_clint_s_xactor_f_rd_data_D_OUT;
  wire soc_clint_s_xactor_f_rd_data_CLR,
       soc_clint_s_xactor_f_rd_data_DEQ,
       soc_clint_s_xactor_f_rd_data_EMPTY_N,
       soc_clint_s_xactor_f_rd_data_ENQ,
       soc_clint_s_xactor_f_rd_data_FULL_N;

  // ports of submodule soc_clint_s_xactor_f_wr_addr
  wire [36 : 0] soc_clint_s_xactor_f_wr_addr_D_IN,
		soc_clint_s_xactor_f_wr_addr_D_OUT;
  wire soc_clint_s_xactor_f_wr_addr_CLR,
       soc_clint_s_xactor_f_wr_addr_DEQ,
       soc_clint_s_xactor_f_wr_addr_EMPTY_N,
       soc_clint_s_xactor_f_wr_addr_ENQ,
       soc_clint_s_xactor_f_wr_addr_FULL_N;

  // ports of submodule soc_clint_s_xactor_f_wr_data
  wire [71 : 0] soc_clint_s_xactor_f_wr_data_D_IN,
		soc_clint_s_xactor_f_wr_data_D_OUT;
  wire soc_clint_s_xactor_f_wr_data_CLR,
       soc_clint_s_xactor_f_wr_data_DEQ,
       soc_clint_s_xactor_f_wr_data_EMPTY_N,
       soc_clint_s_xactor_f_wr_data_ENQ,
       soc_clint_s_xactor_f_wr_data_FULL_N;

  // ports of submodule soc_clint_s_xactor_f_wr_resp
  wire [1 : 0] soc_clint_s_xactor_f_wr_resp_D_IN,
	       soc_clint_s_xactor_f_wr_resp_D_OUT;
  wire soc_clint_s_xactor_f_wr_resp_CLR,
       soc_clint_s_xactor_f_wr_resp_DEQ,
       soc_clint_s_xactor_f_wr_resp_EMPTY_N,
       soc_clint_s_xactor_f_wr_resp_ENQ,
       soc_clint_s_xactor_f_wr_resp_FULL_N;

  // ports of submodule soc_eclass
  wire [63 : 0] soc_eclass_master_d_m_rvalid_rdata,
		soc_eclass_master_d_wdata,
		soc_eclass_master_i_m_rvalid_rdata,
		soc_eclass_master_i_wdata,
		soc_eclass_sb_clint_mtime_put;
  wire [31 : 0] soc_eclass_master_d_araddr,
		soc_eclass_master_d_awaddr,
		soc_eclass_master_i_araddr,
		soc_eclass_master_i_awaddr;
  wire [7 : 0] soc_eclass_master_d_wstrb, soc_eclass_master_i_wstrb;
  wire [2 : 0] soc_eclass_master_d_arprot,
	       soc_eclass_master_d_awprot,
	       soc_eclass_master_i_arprot,
	       soc_eclass_master_i_awprot;
  wire [1 : 0] soc_eclass_master_d_arsize,
	       soc_eclass_master_d_awsize,
	       soc_eclass_master_d_m_bvalid_bresp,
	       soc_eclass_master_d_m_rvalid_rresp,
	       soc_eclass_master_i_arsize,
	       soc_eclass_master_i_awsize,
	       soc_eclass_master_i_m_bvalid_bresp,
	       soc_eclass_master_i_m_rvalid_rresp;
  wire soc_eclass_EN_io_dump_get,
       soc_eclass_EN_sb_clint_msip_put,
       soc_eclass_EN_sb_clint_mtime_put,
       soc_eclass_EN_sb_clint_mtip_put,
       soc_eclass_EN_sb_ext_interrupt_put,
       soc_eclass_master_d_arvalid,
       soc_eclass_master_d_awvalid,
       soc_eclass_master_d_bready,
       soc_eclass_master_d_m_arready_arready,
       soc_eclass_master_d_m_awready_awready,
       soc_eclass_master_d_m_bvalid_bvalid,
       soc_eclass_master_d_m_rvalid_rvalid,
       soc_eclass_master_d_m_wready_wready,
       soc_eclass_master_d_rready,
       soc_eclass_master_d_wvalid,
       soc_eclass_master_i_arvalid,
       soc_eclass_master_i_awvalid,
       soc_eclass_master_i_bready,
       soc_eclass_master_i_m_arready_arready,
       soc_eclass_master_i_m_awready_awready,
       soc_eclass_master_i_m_bvalid_bvalid,
       soc_eclass_master_i_m_rvalid_rvalid,
       soc_eclass_master_i_m_wready_wready,
       soc_eclass_master_i_rready,
       soc_eclass_master_i_wvalid,
       soc_eclass_sb_clint_msip_put,
       soc_eclass_sb_clint_mtip_put,
       soc_eclass_sb_ext_interrupt_put;

  // ports of submodule soc_err_slave_s_xactor_f_rd_addr
  wire [36 : 0] soc_err_slave_s_xactor_f_rd_addr_D_IN;
  wire soc_err_slave_s_xactor_f_rd_addr_CLR,
       soc_err_slave_s_xactor_f_rd_addr_DEQ,
       soc_err_slave_s_xactor_f_rd_addr_EMPTY_N,
       soc_err_slave_s_xactor_f_rd_addr_ENQ,
       soc_err_slave_s_xactor_f_rd_addr_FULL_N;

  // ports of submodule soc_err_slave_s_xactor_f_rd_data
  wire [65 : 0] soc_err_slave_s_xactor_f_rd_data_D_IN,
		soc_err_slave_s_xactor_f_rd_data_D_OUT;
  wire soc_err_slave_s_xactor_f_rd_data_CLR,
       soc_err_slave_s_xactor_f_rd_data_DEQ,
       soc_err_slave_s_xactor_f_rd_data_EMPTY_N,
       soc_err_slave_s_xactor_f_rd_data_ENQ,
       soc_err_slave_s_xactor_f_rd_data_FULL_N;

  // ports of submodule soc_err_slave_s_xactor_f_wr_addr
  wire [36 : 0] soc_err_slave_s_xactor_f_wr_addr_D_IN;
  wire soc_err_slave_s_xactor_f_wr_addr_CLR,
       soc_err_slave_s_xactor_f_wr_addr_DEQ,
       soc_err_slave_s_xactor_f_wr_addr_EMPTY_N,
       soc_err_slave_s_xactor_f_wr_addr_ENQ,
       soc_err_slave_s_xactor_f_wr_addr_FULL_N;

  // ports of submodule soc_err_slave_s_xactor_f_wr_data
  wire [71 : 0] soc_err_slave_s_xactor_f_wr_data_D_IN;
  wire soc_err_slave_s_xactor_f_wr_data_CLR,
       soc_err_slave_s_xactor_f_wr_data_DEQ,
       soc_err_slave_s_xactor_f_wr_data_EMPTY_N,
       soc_err_slave_s_xactor_f_wr_data_ENQ,
       soc_err_slave_s_xactor_f_wr_data_FULL_N;

  // ports of submodule soc_err_slave_s_xactor_f_wr_resp
  wire [1 : 0] soc_err_slave_s_xactor_f_wr_resp_D_IN,
	       soc_err_slave_s_xactor_f_wr_resp_D_OUT;
  wire soc_err_slave_s_xactor_f_wr_resp_CLR,
       soc_err_slave_s_xactor_f_wr_resp_DEQ,
       soc_err_slave_s_xactor_f_wr_resp_EMPTY_N,
       soc_err_slave_s_xactor_f_wr_resp_ENQ,
       soc_err_slave_s_xactor_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_err_user_0
  wire soc_fabric_v_f_rd_err_user_0_CLR,
       soc_fabric_v_f_rd_err_user_0_DEQ,
       soc_fabric_v_f_rd_err_user_0_ENQ;

  // ports of submodule soc_fabric_v_f_rd_err_user_1
  wire soc_fabric_v_f_rd_err_user_1_CLR,
       soc_fabric_v_f_rd_err_user_1_DEQ,
       soc_fabric_v_f_rd_err_user_1_ENQ;

  // ports of submodule soc_fabric_v_f_rd_err_user_2
  wire soc_fabric_v_f_rd_err_user_2_CLR,
       soc_fabric_v_f_rd_err_user_2_DEQ,
       soc_fabric_v_f_rd_err_user_2_ENQ;

  // ports of submodule soc_fabric_v_f_rd_mis_0
  reg [1 : 0] soc_fabric_v_f_rd_mis_0_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_0_D_OUT;
  wire soc_fabric_v_f_rd_mis_0_CLR,
       soc_fabric_v_f_rd_mis_0_DEQ,
       soc_fabric_v_f_rd_mis_0_EMPTY_N,
       soc_fabric_v_f_rd_mis_0_ENQ,
       soc_fabric_v_f_rd_mis_0_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_mis_1
  reg [1 : 0] soc_fabric_v_f_rd_mis_1_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_1_D_OUT;
  wire soc_fabric_v_f_rd_mis_1_CLR,
       soc_fabric_v_f_rd_mis_1_DEQ,
       soc_fabric_v_f_rd_mis_1_EMPTY_N,
       soc_fabric_v_f_rd_mis_1_ENQ,
       soc_fabric_v_f_rd_mis_1_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_mis_2
  reg [1 : 0] soc_fabric_v_f_rd_mis_2_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_2_D_OUT;
  wire soc_fabric_v_f_rd_mis_2_CLR,
       soc_fabric_v_f_rd_mis_2_DEQ,
       soc_fabric_v_f_rd_mis_2_EMPTY_N,
       soc_fabric_v_f_rd_mis_2_ENQ,
       soc_fabric_v_f_rd_mis_2_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_mis_3
  reg [1 : 0] soc_fabric_v_f_rd_mis_3_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_3_D_OUT;
  wire soc_fabric_v_f_rd_mis_3_CLR,
       soc_fabric_v_f_rd_mis_3_DEQ,
       soc_fabric_v_f_rd_mis_3_EMPTY_N,
       soc_fabric_v_f_rd_mis_3_ENQ,
       soc_fabric_v_f_rd_mis_3_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_mis_4
  reg [1 : 0] soc_fabric_v_f_rd_mis_4_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_4_D_OUT;
  wire soc_fabric_v_f_rd_mis_4_CLR,
       soc_fabric_v_f_rd_mis_4_DEQ,
       soc_fabric_v_f_rd_mis_4_EMPTY_N,
       soc_fabric_v_f_rd_mis_4_ENQ,
       soc_fabric_v_f_rd_mis_4_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_mis_5
  reg [1 : 0] soc_fabric_v_f_rd_mis_5_D_IN;
  wire [1 : 0] soc_fabric_v_f_rd_mis_5_D_OUT;
  wire soc_fabric_v_f_rd_mis_5_CLR,
       soc_fabric_v_f_rd_mis_5_DEQ,
       soc_fabric_v_f_rd_mis_5_EMPTY_N,
       soc_fabric_v_f_rd_mis_5_ENQ,
       soc_fabric_v_f_rd_mis_5_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_sjs_0
  reg [2 : 0] soc_fabric_v_f_rd_sjs_0_D_IN;
  wire [2 : 0] soc_fabric_v_f_rd_sjs_0_D_OUT;
  wire soc_fabric_v_f_rd_sjs_0_CLR,
       soc_fabric_v_f_rd_sjs_0_DEQ,
       soc_fabric_v_f_rd_sjs_0_EMPTY_N,
       soc_fabric_v_f_rd_sjs_0_ENQ,
       soc_fabric_v_f_rd_sjs_0_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_sjs_1
  reg [2 : 0] soc_fabric_v_f_rd_sjs_1_D_IN;
  wire [2 : 0] soc_fabric_v_f_rd_sjs_1_D_OUT;
  wire soc_fabric_v_f_rd_sjs_1_CLR,
       soc_fabric_v_f_rd_sjs_1_DEQ,
       soc_fabric_v_f_rd_sjs_1_EMPTY_N,
       soc_fabric_v_f_rd_sjs_1_ENQ,
       soc_fabric_v_f_rd_sjs_1_FULL_N;

  // ports of submodule soc_fabric_v_f_rd_sjs_2
  reg [2 : 0] soc_fabric_v_f_rd_sjs_2_D_IN;
  wire [2 : 0] soc_fabric_v_f_rd_sjs_2_D_OUT;
  wire soc_fabric_v_f_rd_sjs_2_CLR,
       soc_fabric_v_f_rd_sjs_2_DEQ,
       soc_fabric_v_f_rd_sjs_2_EMPTY_N,
       soc_fabric_v_f_rd_sjs_2_ENQ,
       soc_fabric_v_f_rd_sjs_2_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_err_user_0
  wire soc_fabric_v_f_wr_err_user_0_CLR,
       soc_fabric_v_f_wr_err_user_0_DEQ,
       soc_fabric_v_f_wr_err_user_0_ENQ;

  // ports of submodule soc_fabric_v_f_wr_err_user_1
  wire soc_fabric_v_f_wr_err_user_1_CLR,
       soc_fabric_v_f_wr_err_user_1_DEQ,
       soc_fabric_v_f_wr_err_user_1_ENQ;

  // ports of submodule soc_fabric_v_f_wr_err_user_2
  wire soc_fabric_v_f_wr_err_user_2_CLR,
       soc_fabric_v_f_wr_err_user_2_DEQ,
       soc_fabric_v_f_wr_err_user_2_ENQ;

  // ports of submodule soc_fabric_v_f_wr_mis_0
  reg [1 : 0] soc_fabric_v_f_wr_mis_0_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_0_D_OUT;
  wire soc_fabric_v_f_wr_mis_0_CLR,
       soc_fabric_v_f_wr_mis_0_DEQ,
       soc_fabric_v_f_wr_mis_0_EMPTY_N,
       soc_fabric_v_f_wr_mis_0_ENQ,
       soc_fabric_v_f_wr_mis_0_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_mis_1
  reg [1 : 0] soc_fabric_v_f_wr_mis_1_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_1_D_OUT;
  wire soc_fabric_v_f_wr_mis_1_CLR,
       soc_fabric_v_f_wr_mis_1_DEQ,
       soc_fabric_v_f_wr_mis_1_EMPTY_N,
       soc_fabric_v_f_wr_mis_1_ENQ,
       soc_fabric_v_f_wr_mis_1_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_mis_2
  reg [1 : 0] soc_fabric_v_f_wr_mis_2_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_2_D_OUT;
  wire soc_fabric_v_f_wr_mis_2_CLR,
       soc_fabric_v_f_wr_mis_2_DEQ,
       soc_fabric_v_f_wr_mis_2_EMPTY_N,
       soc_fabric_v_f_wr_mis_2_ENQ,
       soc_fabric_v_f_wr_mis_2_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_mis_3
  reg [1 : 0] soc_fabric_v_f_wr_mis_3_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_3_D_OUT;
  wire soc_fabric_v_f_wr_mis_3_CLR,
       soc_fabric_v_f_wr_mis_3_DEQ,
       soc_fabric_v_f_wr_mis_3_EMPTY_N,
       soc_fabric_v_f_wr_mis_3_ENQ,
       soc_fabric_v_f_wr_mis_3_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_mis_4
  reg [1 : 0] soc_fabric_v_f_wr_mis_4_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_4_D_OUT;
  wire soc_fabric_v_f_wr_mis_4_CLR,
       soc_fabric_v_f_wr_mis_4_DEQ,
       soc_fabric_v_f_wr_mis_4_EMPTY_N,
       soc_fabric_v_f_wr_mis_4_ENQ,
       soc_fabric_v_f_wr_mis_4_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_mis_5
  reg [1 : 0] soc_fabric_v_f_wr_mis_5_D_IN;
  wire [1 : 0] soc_fabric_v_f_wr_mis_5_D_OUT;
  wire soc_fabric_v_f_wr_mis_5_CLR,
       soc_fabric_v_f_wr_mis_5_DEQ,
       soc_fabric_v_f_wr_mis_5_EMPTY_N,
       soc_fabric_v_f_wr_mis_5_ENQ,
       soc_fabric_v_f_wr_mis_5_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_sjs_0
  reg [2 : 0] soc_fabric_v_f_wr_sjs_0_D_IN;
  wire [2 : 0] soc_fabric_v_f_wr_sjs_0_D_OUT;
  wire soc_fabric_v_f_wr_sjs_0_CLR,
       soc_fabric_v_f_wr_sjs_0_DEQ,
       soc_fabric_v_f_wr_sjs_0_EMPTY_N,
       soc_fabric_v_f_wr_sjs_0_ENQ,
       soc_fabric_v_f_wr_sjs_0_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_sjs_1
  reg [2 : 0] soc_fabric_v_f_wr_sjs_1_D_IN;
  wire [2 : 0] soc_fabric_v_f_wr_sjs_1_D_OUT;
  wire soc_fabric_v_f_wr_sjs_1_CLR,
       soc_fabric_v_f_wr_sjs_1_DEQ,
       soc_fabric_v_f_wr_sjs_1_EMPTY_N,
       soc_fabric_v_f_wr_sjs_1_ENQ,
       soc_fabric_v_f_wr_sjs_1_FULL_N;

  // ports of submodule soc_fabric_v_f_wr_sjs_2
  reg [2 : 0] soc_fabric_v_f_wr_sjs_2_D_IN;
  wire [2 : 0] soc_fabric_v_f_wr_sjs_2_D_OUT;
  wire soc_fabric_v_f_wr_sjs_2_CLR,
       soc_fabric_v_f_wr_sjs_2_DEQ,
       soc_fabric_v_f_wr_sjs_2_EMPTY_N,
       soc_fabric_v_f_wr_sjs_2_ENQ,
       soc_fabric_v_f_wr_sjs_2_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_0_f_rd_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_0_f_rd_addr_D_IN,
		soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_0_f_rd_addr_CLR,
       soc_fabric_xactors_from_masters_0_f_rd_addr_DEQ,
       soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_0_f_rd_addr_ENQ,
       soc_fabric_xactors_from_masters_0_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_0_f_rd_data
  reg [65 : 0] soc_fabric_xactors_from_masters_0_f_rd_data_D_IN;
  wire [65 : 0] soc_fabric_xactors_from_masters_0_f_rd_data_D_OUT;
  wire soc_fabric_xactors_from_masters_0_f_rd_data_CLR,
       soc_fabric_xactors_from_masters_0_f_rd_data_DEQ,
       soc_fabric_xactors_from_masters_0_f_rd_data_EMPTY_N,
       soc_fabric_xactors_from_masters_0_f_rd_data_ENQ,
       soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_0_f_wr_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_0_f_wr_addr_D_IN,
		soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_0_f_wr_addr_CLR,
       soc_fabric_xactors_from_masters_0_f_wr_addr_DEQ,
       soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_0_f_wr_addr_ENQ,
       soc_fabric_xactors_from_masters_0_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_0_f_wr_data
  wire [71 : 0] soc_fabric_xactors_from_masters_0_f_wr_data_D_IN,
		soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
  wire soc_fabric_xactors_from_masters_0_f_wr_data_CLR,
       soc_fabric_xactors_from_masters_0_f_wr_data_DEQ,
       soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N,
       soc_fabric_xactors_from_masters_0_f_wr_data_ENQ,
       soc_fabric_xactors_from_masters_0_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_0_f_wr_resp
  reg [1 : 0] soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN;
  wire [1 : 0] soc_fabric_xactors_from_masters_0_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_from_masters_0_f_wr_resp_CLR,
       soc_fabric_xactors_from_masters_0_f_wr_resp_DEQ,
       soc_fabric_xactors_from_masters_0_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_from_masters_0_f_wr_resp_ENQ,
       soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_1_f_rd_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_1_f_rd_addr_D_IN,
		soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_1_f_rd_addr_CLR,
       soc_fabric_xactors_from_masters_1_f_rd_addr_DEQ,
       soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_1_f_rd_addr_ENQ,
       soc_fabric_xactors_from_masters_1_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_1_f_rd_data
  reg [65 : 0] soc_fabric_xactors_from_masters_1_f_rd_data_D_IN;
  wire [65 : 0] soc_fabric_xactors_from_masters_1_f_rd_data_D_OUT;
  wire soc_fabric_xactors_from_masters_1_f_rd_data_CLR,
       soc_fabric_xactors_from_masters_1_f_rd_data_DEQ,
       soc_fabric_xactors_from_masters_1_f_rd_data_EMPTY_N,
       soc_fabric_xactors_from_masters_1_f_rd_data_ENQ,
       soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_1_f_wr_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_1_f_wr_addr_D_IN,
		soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_1_f_wr_addr_CLR,
       soc_fabric_xactors_from_masters_1_f_wr_addr_DEQ,
       soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_1_f_wr_addr_ENQ,
       soc_fabric_xactors_from_masters_1_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_1_f_wr_data
  wire [71 : 0] soc_fabric_xactors_from_masters_1_f_wr_data_D_IN,
		soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
  wire soc_fabric_xactors_from_masters_1_f_wr_data_CLR,
       soc_fabric_xactors_from_masters_1_f_wr_data_DEQ,
       soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N,
       soc_fabric_xactors_from_masters_1_f_wr_data_ENQ,
       soc_fabric_xactors_from_masters_1_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_1_f_wr_resp
  reg [1 : 0] soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN;
  wire [1 : 0] soc_fabric_xactors_from_masters_1_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_from_masters_1_f_wr_resp_CLR,
       soc_fabric_xactors_from_masters_1_f_wr_resp_DEQ,
       soc_fabric_xactors_from_masters_1_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_from_masters_1_f_wr_resp_ENQ,
       soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_2_f_rd_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_2_f_rd_addr_D_IN,
		soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_2_f_rd_addr_CLR,
       soc_fabric_xactors_from_masters_2_f_rd_addr_DEQ,
       soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_2_f_rd_addr_ENQ,
       soc_fabric_xactors_from_masters_2_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_2_f_rd_data
  reg [65 : 0] soc_fabric_xactors_from_masters_2_f_rd_data_D_IN;
  wire [65 : 0] soc_fabric_xactors_from_masters_2_f_rd_data_D_OUT;
  wire soc_fabric_xactors_from_masters_2_f_rd_data_CLR,
       soc_fabric_xactors_from_masters_2_f_rd_data_DEQ,
       soc_fabric_xactors_from_masters_2_f_rd_data_EMPTY_N,
       soc_fabric_xactors_from_masters_2_f_rd_data_ENQ,
       soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_2_f_wr_addr
  wire [36 : 0] soc_fabric_xactors_from_masters_2_f_wr_addr_D_IN,
		soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_from_masters_2_f_wr_addr_CLR,
       soc_fabric_xactors_from_masters_2_f_wr_addr_DEQ,
       soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_from_masters_2_f_wr_addr_ENQ,
       soc_fabric_xactors_from_masters_2_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_2_f_wr_data
  wire [71 : 0] soc_fabric_xactors_from_masters_2_f_wr_data_D_IN,
		soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
  wire soc_fabric_xactors_from_masters_2_f_wr_data_CLR,
       soc_fabric_xactors_from_masters_2_f_wr_data_DEQ,
       soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N,
       soc_fabric_xactors_from_masters_2_f_wr_data_ENQ,
       soc_fabric_xactors_from_masters_2_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_from_masters_2_f_wr_resp
  reg [1 : 0] soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN;
  wire [1 : 0] soc_fabric_xactors_from_masters_2_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_from_masters_2_f_wr_resp_CLR,
       soc_fabric_xactors_from_masters_2_f_wr_resp_DEQ,
       soc_fabric_xactors_from_masters_2_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_from_masters_2_f_wr_resp_ENQ,
       soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_0_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN;
  wire soc_fabric_xactors_to_slaves_0_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_0_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_0_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_0_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_0_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_0_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_0_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_0_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_0_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_0_f_rd_data_ENQ;

  // ports of submodule soc_fabric_xactors_to_slaves_0_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN;
  wire soc_fabric_xactors_to_slaves_0_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_0_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_0_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_0_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_0_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN;
  wire soc_fabric_xactors_to_slaves_0_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_0_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_0_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_0_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_0_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_0_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_0_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_0_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_0_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_0_f_wr_resp_ENQ;

  // ports of submodule soc_fabric_xactors_to_slaves_1_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN;
  wire soc_fabric_xactors_to_slaves_1_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_1_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_1_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_1_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_1_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_1_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_1_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_1_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_1_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_1_f_rd_data_ENQ;

  // ports of submodule soc_fabric_xactors_to_slaves_1_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN;
  wire soc_fabric_xactors_to_slaves_1_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_1_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_1_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_1_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_1_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN;
  wire soc_fabric_xactors_to_slaves_1_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_1_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_1_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_1_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_1_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_1_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_1_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_1_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_1_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_1_f_wr_resp_ENQ;

  // ports of submodule soc_fabric_xactors_to_slaves_2_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_2_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_2_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_2_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_2_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_2_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_2_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_2_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_2_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_2_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_2_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_2_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_2_f_rd_data_ENQ,
       soc_fabric_xactors_to_slaves_2_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_2_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_2_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_2_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_2_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_2_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_2_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_2_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_2_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN;
  wire [71 : 0] soc_fabric_xactors_to_slaves_2_f_wr_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_2_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_2_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_2_f_wr_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_2_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_2_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_2_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_2_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_2_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_2_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_2_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_2_f_wr_resp_ENQ,
       soc_fabric_xactors_to_slaves_2_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_3_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_3_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_3_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_3_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_3_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_3_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_3_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_3_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_3_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_3_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_3_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_3_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_3_f_rd_data_ENQ,
       soc_fabric_xactors_to_slaves_3_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_3_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_3_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_3_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_3_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_3_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_3_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_3_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_3_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN;
  wire [71 : 0] soc_fabric_xactors_to_slaves_3_f_wr_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_3_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_3_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_3_f_wr_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_3_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_3_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_3_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_3_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_3_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_3_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_3_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_3_f_wr_resp_ENQ,
       soc_fabric_xactors_to_slaves_3_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_4_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_4_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_4_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_4_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_4_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_4_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_4_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_4_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_4_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_4_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_4_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_4_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_4_f_rd_data_ENQ,
       soc_fabric_xactors_to_slaves_4_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_4_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_4_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_4_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_4_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_4_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_4_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_4_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_4_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN;
  wire [71 : 0] soc_fabric_xactors_to_slaves_4_f_wr_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_4_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_4_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_4_f_wr_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_4_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_4_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_4_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_4_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_4_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_4_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_4_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_4_f_wr_resp_ENQ,
       soc_fabric_xactors_to_slaves_4_f_wr_resp_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_5_f_rd_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_5_f_rd_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_5_f_rd_addr_CLR,
       soc_fabric_xactors_to_slaves_5_f_rd_addr_DEQ,
       soc_fabric_xactors_to_slaves_5_f_rd_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_5_f_rd_addr_ENQ,
       soc_fabric_xactors_to_slaves_5_f_rd_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_5_f_rd_data
  wire [65 : 0] soc_fabric_xactors_to_slaves_5_f_rd_data_D_IN,
		soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_5_f_rd_data_CLR,
       soc_fabric_xactors_to_slaves_5_f_rd_data_DEQ,
       soc_fabric_xactors_to_slaves_5_f_rd_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_5_f_rd_data_ENQ,
       soc_fabric_xactors_to_slaves_5_f_rd_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_5_f_wr_addr
  reg [36 : 0] soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN;
  wire [36 : 0] soc_fabric_xactors_to_slaves_5_f_wr_addr_D_OUT;
  wire soc_fabric_xactors_to_slaves_5_f_wr_addr_CLR,
       soc_fabric_xactors_to_slaves_5_f_wr_addr_DEQ,
       soc_fabric_xactors_to_slaves_5_f_wr_addr_EMPTY_N,
       soc_fabric_xactors_to_slaves_5_f_wr_addr_ENQ,
       soc_fabric_xactors_to_slaves_5_f_wr_addr_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_5_f_wr_data
  reg [71 : 0] soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN;
  wire [71 : 0] soc_fabric_xactors_to_slaves_5_f_wr_data_D_OUT;
  wire soc_fabric_xactors_to_slaves_5_f_wr_data_CLR,
       soc_fabric_xactors_to_slaves_5_f_wr_data_DEQ,
       soc_fabric_xactors_to_slaves_5_f_wr_data_EMPTY_N,
       soc_fabric_xactors_to_slaves_5_f_wr_data_ENQ,
       soc_fabric_xactors_to_slaves_5_f_wr_data_FULL_N;

  // ports of submodule soc_fabric_xactors_to_slaves_5_f_wr_resp
  wire [1 : 0] soc_fabric_xactors_to_slaves_5_f_wr_resp_D_IN,
	       soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT;
  wire soc_fabric_xactors_to_slaves_5_f_wr_resp_CLR,
       soc_fabric_xactors_to_slaves_5_f_wr_resp_DEQ,
       soc_fabric_xactors_to_slaves_5_f_wr_resp_EMPTY_N,
       soc_fabric_xactors_to_slaves_5_f_wr_resp_ENQ,
       soc_fabric_xactors_to_slaves_5_f_wr_resp_FULL_N;

  // ports of submodule soc_signature
  wire [63 : 0] soc_signature_master_m_rvalid_rdata,
		soc_signature_master_wdata,
		soc_signature_slave_m_wvalid_wdata,
		soc_signature_slave_rdata;
  wire [31 : 0] soc_signature_master_araddr,
		soc_signature_master_awaddr,
		soc_signature_slave_m_arvalid_araddr,
		soc_signature_slave_m_awvalid_awaddr;
  wire [7 : 0] soc_signature_master_wstrb, soc_signature_slave_m_wvalid_wstrb;
  wire [2 : 0] soc_signature_master_arprot,
	       soc_signature_master_awprot,
	       soc_signature_slave_m_arvalid_arprot,
	       soc_signature_slave_m_awvalid_awprot;
  wire [1 : 0] soc_signature_master_arsize,
	       soc_signature_master_awsize,
	       soc_signature_master_m_bvalid_bresp,
	       soc_signature_master_m_rvalid_rresp,
	       soc_signature_slave_bresp,
	       soc_signature_slave_m_arvalid_arsize,
	       soc_signature_slave_m_awvalid_awsize,
	       soc_signature_slave_rresp;
  wire soc_signature_master_arvalid,
       soc_signature_master_awvalid,
       soc_signature_master_bready,
       soc_signature_master_m_arready_arready,
       soc_signature_master_m_awready_awready,
       soc_signature_master_m_bvalid_bvalid,
       soc_signature_master_m_rvalid_rvalid,
       soc_signature_master_m_wready_wready,
       soc_signature_master_rready,
       soc_signature_master_wvalid,
       soc_signature_slave_arready,
       soc_signature_slave_awready,
       soc_signature_slave_bvalid,
       soc_signature_slave_m_arvalid_arvalid,
       soc_signature_slave_m_awvalid_awvalid,
       soc_signature_slave_m_bready_bready,
       soc_signature_slave_m_rready_rready,
       soc_signature_slave_m_wvalid_wvalid,
       soc_signature_slave_rvalid,
       soc_signature_slave_wready;

  // ports of submodule soc_uart_s_xactor_f_rd_addr
  wire [36 : 0] soc_uart_s_xactor_f_rd_addr_D_IN,
		soc_uart_s_xactor_f_rd_addr_D_OUT;
  wire soc_uart_s_xactor_f_rd_addr_CLR,
       soc_uart_s_xactor_f_rd_addr_DEQ,
       soc_uart_s_xactor_f_rd_addr_EMPTY_N,
       soc_uart_s_xactor_f_rd_addr_ENQ,
       soc_uart_s_xactor_f_rd_addr_FULL_N;

  // ports of submodule soc_uart_s_xactor_f_rd_data
  wire [65 : 0] soc_uart_s_xactor_f_rd_data_D_IN,
		soc_uart_s_xactor_f_rd_data_D_OUT;
  wire soc_uart_s_xactor_f_rd_data_CLR,
       soc_uart_s_xactor_f_rd_data_DEQ,
       soc_uart_s_xactor_f_rd_data_EMPTY_N,
       soc_uart_s_xactor_f_rd_data_ENQ,
       soc_uart_s_xactor_f_rd_data_FULL_N;

  // ports of submodule soc_uart_s_xactor_f_wr_addr
  wire [36 : 0] soc_uart_s_xactor_f_wr_addr_D_IN,
		soc_uart_s_xactor_f_wr_addr_D_OUT;
  wire soc_uart_s_xactor_f_wr_addr_CLR,
       soc_uart_s_xactor_f_wr_addr_DEQ,
       soc_uart_s_xactor_f_wr_addr_EMPTY_N,
       soc_uart_s_xactor_f_wr_addr_ENQ,
       soc_uart_s_xactor_f_wr_addr_FULL_N;

  // ports of submodule soc_uart_s_xactor_f_wr_data
  wire [71 : 0] soc_uart_s_xactor_f_wr_data_D_IN,
		soc_uart_s_xactor_f_wr_data_D_OUT;
  wire soc_uart_s_xactor_f_wr_data_CLR,
       soc_uart_s_xactor_f_wr_data_DEQ,
       soc_uart_s_xactor_f_wr_data_EMPTY_N,
       soc_uart_s_xactor_f_wr_data_ENQ,
       soc_uart_s_xactor_f_wr_data_FULL_N;

  // ports of submodule soc_uart_s_xactor_f_wr_resp
  wire [1 : 0] soc_uart_s_xactor_f_wr_resp_D_IN,
	       soc_uart_s_xactor_f_wr_resp_D_OUT;
  wire soc_uart_s_xactor_f_wr_resp_CLR,
       soc_uart_s_xactor_f_wr_resp_DEQ,
       soc_uart_s_xactor_f_wr_resp_EMPTY_N,
       soc_uart_s_xactor_f_wr_resp_ENQ,
       soc_uart_s_xactor_f_wr_resp_FULL_N;

  // ports of submodule soc_uart_user_ifc_uart_baudGen_rBaudCounter
  wire [15 : 0] soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_A,
		soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_B,
		soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_C,
		soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_F,
		soc_uart_user_ifc_uart_baudGen_rBaudCounter_Q_OUT;
  wire soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDA,
       soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDB,
       soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETC,
       soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETF;

  // ports of submodule soc_uart_user_ifc_uart_baudGen_rBaudTickCounter
  wire [2 : 0] soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_A,
	       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_B,
	       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_C,
	       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_F,
	       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_Q_OUT;
  wire soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDA,
       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDB,
       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETC,
       soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETF;

  // ports of submodule soc_uart_user_ifc_uart_fifoRecv
  wire [7 : 0] soc_uart_user_ifc_uart_fifoRecv_D_IN,
	       soc_uart_user_ifc_uart_fifoRecv_D_OUT;
  wire soc_uart_user_ifc_uart_fifoRecv_CLR,
       soc_uart_user_ifc_uart_fifoRecv_DEQ,
       soc_uart_user_ifc_uart_fifoRecv_EMPTY_N,
       soc_uart_user_ifc_uart_fifoRecv_ENQ,
       soc_uart_user_ifc_uart_fifoRecv_FULL_N;

  // ports of submodule soc_uart_user_ifc_uart_fifoXmit
  wire [7 : 0] soc_uart_user_ifc_uart_fifoXmit_D_IN,
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT;
  wire soc_uart_user_ifc_uart_fifoXmit_CLR,
       soc_uart_user_ifc_uart_fifoXmit_DEQ,
       soc_uart_user_ifc_uart_fifoXmit_EMPTY_N,
       soc_uart_user_ifc_uart_fifoXmit_ENQ,
       soc_uart_user_ifc_uart_fifoXmit_FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_soc_1_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_1_rl_rd_data_channel,
       CAN_FIRE_RL_soc_1_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_1_rl_wr_data_channel,
       CAN_FIRE_RL_soc_1_rl_wr_response_channel,
       CAN_FIRE_RL_soc_2_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_2_rl_rd_data_channel,
       CAN_FIRE_RL_soc_2_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_2_rl_wr_data_channel,
       CAN_FIRE_RL_soc_2_rl_wr_response_channel,
       CAN_FIRE_RL_soc_3_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_3_rl_rd_data_channel,
       CAN_FIRE_RL_soc_3_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_3_rl_wr_data_channel,
       CAN_FIRE_RL_soc_3_rl_wr_response_channel,
       CAN_FIRE_RL_soc_4_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_4_rl_rd_data_channel,
       CAN_FIRE_RL_soc_4_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_4_rl_wr_data_channel,
       CAN_FIRE_RL_soc_4_rl_wr_response_channel,
       CAN_FIRE_RL_soc_5_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_5_rl_rd_data_channel,
       CAN_FIRE_RL_soc_5_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_5_rl_wr_data_channel,
       CAN_FIRE_RL_soc_5_rl_wr_response_channel,
       CAN_FIRE_RL_soc_6_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_6_rl_rd_data_channel,
       CAN_FIRE_RL_soc_6_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_6_rl_wr_data_channel,
       CAN_FIRE_RL_soc_6_rl_wr_response_channel,
       CAN_FIRE_RL_soc_7_mkConnectionGetPut,
       CAN_FIRE_RL_soc_8_mkConnectionGetPut,
       CAN_FIRE_RL_soc_9_mkConnectionGetPut,
       CAN_FIRE_RL_soc_clint_axi_read_transaction,
       CAN_FIRE_RL_soc_clint_axi_write_transaction,
       CAN_FIRE_RL_soc_clint_clint_clear_interrupt,
       CAN_FIRE_RL_soc_clint_clint_generate_time_interrupt,
       CAN_FIRE_RL_soc_clint_clint_increment_timer,
       CAN_FIRE_RL_soc_err_slave_receive_read_request,
       CAN_FIRE_RL_soc_err_slave_receive_write_request,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8,
       CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8,
       CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8,
       CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8,
       CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9,
       CAN_FIRE_RL_soc_rl_rd_addr_channel,
       CAN_FIRE_RL_soc_rl_rd_data_channel,
       CAN_FIRE_RL_soc_rl_wr_addr_channel,
       CAN_FIRE_RL_soc_rl_wr_data_channel,
       CAN_FIRE_RL_soc_rl_wr_response_channel,
       CAN_FIRE_RL_soc_uart_capture_read_request,
       CAN_FIRE_RL_soc_uart_capture_write_request,
       CAN_FIRE_RL_soc_uart_user_ifc_capture_status,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_count_wire,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_tick_count_wire,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_baud_generator_clock_enable,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_cell_time_counter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_counter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_cell_time_counter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_counter,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time,
       CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command,
       WILL_FIRE_RL_soc_1_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_1_rl_rd_data_channel,
       WILL_FIRE_RL_soc_1_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_1_rl_wr_data_channel,
       WILL_FIRE_RL_soc_1_rl_wr_response_channel,
       WILL_FIRE_RL_soc_2_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_2_rl_rd_data_channel,
       WILL_FIRE_RL_soc_2_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_2_rl_wr_data_channel,
       WILL_FIRE_RL_soc_2_rl_wr_response_channel,
       WILL_FIRE_RL_soc_3_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_3_rl_rd_data_channel,
       WILL_FIRE_RL_soc_3_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_3_rl_wr_data_channel,
       WILL_FIRE_RL_soc_3_rl_wr_response_channel,
       WILL_FIRE_RL_soc_4_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_4_rl_rd_data_channel,
       WILL_FIRE_RL_soc_4_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_4_rl_wr_data_channel,
       WILL_FIRE_RL_soc_4_rl_wr_response_channel,
       WILL_FIRE_RL_soc_5_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_5_rl_rd_data_channel,
       WILL_FIRE_RL_soc_5_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_5_rl_wr_data_channel,
       WILL_FIRE_RL_soc_5_rl_wr_response_channel,
       WILL_FIRE_RL_soc_6_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_6_rl_rd_data_channel,
       WILL_FIRE_RL_soc_6_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_6_rl_wr_data_channel,
       WILL_FIRE_RL_soc_6_rl_wr_response_channel,
       WILL_FIRE_RL_soc_7_mkConnectionGetPut,
       WILL_FIRE_RL_soc_8_mkConnectionGetPut,
       WILL_FIRE_RL_soc_9_mkConnectionGetPut,
       WILL_FIRE_RL_soc_clint_axi_read_transaction,
       WILL_FIRE_RL_soc_clint_axi_write_transaction,
       WILL_FIRE_RL_soc_clint_clint_clear_interrupt,
       WILL_FIRE_RL_soc_clint_clint_generate_time_interrupt,
       WILL_FIRE_RL_soc_clint_clint_increment_timer,
       WILL_FIRE_RL_soc_err_slave_receive_read_request,
       WILL_FIRE_RL_soc_err_slave_receive_write_request,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8,
       WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8,
       WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8,
       WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8,
       WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9,
       WILL_FIRE_RL_soc_rl_rd_addr_channel,
       WILL_FIRE_RL_soc_rl_rd_data_channel,
       WILL_FIRE_RL_soc_rl_wr_addr_channel,
       WILL_FIRE_RL_soc_rl_wr_data_channel,
       WILL_FIRE_RL_soc_rl_wr_response_channel,
       WILL_FIRE_RL_soc_uart_capture_read_request,
       WILL_FIRE_RL_soc_uart_capture_write_request,
       WILL_FIRE_RL_soc_uart_user_ifc_capture_status,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_count_wire,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_tick_count_wire,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_baud_generator_clock_enable,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_cell_time_counter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_counter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_cell_time_counter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_counter,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time,
       WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command;

  // inputs to muxes for submodule ports
  reg [2 : 0] MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_3;
  wire [2 : 0] MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_1,
	       MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_2,
	       MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_4,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_1,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_2,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_3,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_4,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_5,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_6,
	       MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_7;
  wire MUX_soc_clint_clint_mtip_write_1__VAL_1,
       MUX_soc_uart_user_ifc_uart_rRecvState_write_1__SEL_6,
       MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_1,
       MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_2,
       MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_3;

  // remaining internal signals
  reg [63 : 0] IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078,
	       data__h56748,
	       mask__h56747;
  wire [63 : 0] IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1070,
		IF_soc_uart_s_xactor_f_rd_addr_first__39_BITS__ETC___d971,
		_theResult___snd__h46661,
		_theResult___snd__h46728,
		_theResult___snd__h46795,
		a__h41688,
		a__h41694,
		a__h41696,
		datamask__h56751,
		mask__h56750,
		notmask__h56752,
		temp___1__h46656,
		temp___1__h47250,
		temp__h46605,
		temp__h46821,
		temp__h56130,
		x__h58828;
  wire [5 : 0] shift_amt__h46602, shift_amt__h56749;
  wire [3 : 0] x__h33749, x__h35390, x__h37182, x__h37208;
  wire _dor2soc_uart_user_ifc_uart_pwXmitCellCountReset_EN_wset,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d296,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d305,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d307,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d310,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d320,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d322,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d325,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d327,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d337,
       soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d339,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d101,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d103,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d51,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d63,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d65,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d68,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d81,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d83,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d86,
       soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d88,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d372,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d378,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d380,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d383,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d390,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d392,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d395,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d397,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d404,
       soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d406,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d142,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d149,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d151,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d154,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d162,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d164,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d167,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d169,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d177,
       soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d179,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d439,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d445,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d447,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d450,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d457,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d459,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d462,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d464,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d471,
       soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d473,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d218,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d225,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d227,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d230,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d238,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d240,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d243,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d245,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d253,
       soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d255,
       soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802,
       z__h38596,
       z__h38603,
       z__h38610,
       z__h38617,
       z__h38624,
       z__h38631;

  // value method rvfi_valid
  assign rvfi_valid = 1'd1 ;

  // value method rvfi_order
  assign rvfi_order = 64'd0 ;

  // value method rvfi_insn
  assign rvfi_insn = 32'd0 ;

  // value method rvfi_trap
  assign rvfi_trap = 1'd0 ;

  // value method rvfi_halt
  assign rvfi_halt = 1'd0 ;

  // value method rvfi_intr
  assign rvfi_intr = 1'd0 ;

  // value method rvfi_mode
  assign rvfi_mode = 2'd3 ;

  // value method rvfi_ixl
  assign rvfi_ixl = 2'd1 ;

  // value method rvfi_mem_addr
  assign rvfi_mem_addr = 32'd0 ;

  // value method rvfi_mem_rmask
  assign rvfi_mem_rmask = 4'd0 ;

  // value method rvfi_mem_wmask
  assign rvfi_mem_wmask = 4'd0 ;

  // value method rvfi_mem_rdata
  assign rvfi_mem_rdata = 32'd0 ;

  // value method rvfi_mem_wdata
  assign rvfi_mem_wdata = 32'd0 ;

  // value method rvfi_rs1_addr
  assign rvfi_rs1_addr = 5'd0 ;

  // value method rvfi_rs2_addr
  assign rvfi_rs2_addr = 5'd0 ;

  // value method rvfi_rs1_rdata
  assign rvfi_rs1_rdata = 32'd0 ;

  // value method rvfi_rs2_rdata
  assign rvfi_rs2_rdata = 32'd0 ;

  // value method rvfi_rd_addr
  assign rvfi_rd_addr = 5'd0 ;

  // value method rvfi_rd_wdata
  assign rvfi_rd_wdata = 32'd0 ;

  // value method rvfi_pc_rdata
  assign rvfi_pc_rdata = 32'd0 ;

  // value method rvfi_pc_wdata
  assign rvfi_pc_wdata = 32'd0 ;

  // submodule soc_clint_s_xactor_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_clint_s_xactor_f_rd_addr(.RST(RST_N),
							.CLK(CLK),
							.D_IN(soc_clint_s_xactor_f_rd_addr_D_IN),
							.ENQ(soc_clint_s_xactor_f_rd_addr_ENQ),
							.DEQ(soc_clint_s_xactor_f_rd_addr_DEQ),
							.CLR(soc_clint_s_xactor_f_rd_addr_CLR),
							.D_OUT(soc_clint_s_xactor_f_rd_addr_D_OUT),
							.FULL_N(soc_clint_s_xactor_f_rd_addr_FULL_N),
							.EMPTY_N(soc_clint_s_xactor_f_rd_addr_EMPTY_N));

  // submodule soc_clint_s_xactor_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_clint_s_xactor_f_rd_data(.RST(RST_N),
							.CLK(CLK),
							.D_IN(soc_clint_s_xactor_f_rd_data_D_IN),
							.ENQ(soc_clint_s_xactor_f_rd_data_ENQ),
							.DEQ(soc_clint_s_xactor_f_rd_data_DEQ),
							.CLR(soc_clint_s_xactor_f_rd_data_CLR),
							.D_OUT(soc_clint_s_xactor_f_rd_data_D_OUT),
							.FULL_N(soc_clint_s_xactor_f_rd_data_FULL_N),
							.EMPTY_N(soc_clint_s_xactor_f_rd_data_EMPTY_N));

  // submodule soc_clint_s_xactor_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_clint_s_xactor_f_wr_addr(.RST(RST_N),
							.CLK(CLK),
							.D_IN(soc_clint_s_xactor_f_wr_addr_D_IN),
							.ENQ(soc_clint_s_xactor_f_wr_addr_ENQ),
							.DEQ(soc_clint_s_xactor_f_wr_addr_DEQ),
							.CLR(soc_clint_s_xactor_f_wr_addr_CLR),
							.D_OUT(soc_clint_s_xactor_f_wr_addr_D_OUT),
							.FULL_N(soc_clint_s_xactor_f_wr_addr_FULL_N),
							.EMPTY_N(soc_clint_s_xactor_f_wr_addr_EMPTY_N));

  // submodule soc_clint_s_xactor_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_clint_s_xactor_f_wr_data(.RST(RST_N),
							.CLK(CLK),
							.D_IN(soc_clint_s_xactor_f_wr_data_D_IN),
							.ENQ(soc_clint_s_xactor_f_wr_data_ENQ),
							.DEQ(soc_clint_s_xactor_f_wr_data_DEQ),
							.CLR(soc_clint_s_xactor_f_wr_data_CLR),
							.D_OUT(soc_clint_s_xactor_f_wr_data_D_OUT),
							.FULL_N(soc_clint_s_xactor_f_wr_data_FULL_N),
							.EMPTY_N(soc_clint_s_xactor_f_wr_data_EMPTY_N));

  // submodule soc_clint_s_xactor_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_clint_s_xactor_f_wr_resp(.RST(RST_N),
							.CLK(CLK),
							.D_IN(soc_clint_s_xactor_f_wr_resp_D_IN),
							.ENQ(soc_clint_s_xactor_f_wr_resp_ENQ),
							.DEQ(soc_clint_s_xactor_f_wr_resp_DEQ),
							.CLR(soc_clint_s_xactor_f_wr_resp_CLR),
							.D_OUT(soc_clint_s_xactor_f_wr_resp_D_OUT),
							.FULL_N(soc_clint_s_xactor_f_wr_resp_FULL_N),
							.EMPTY_N(soc_clint_s_xactor_f_wr_resp_EMPTY_N));

  // submodule soc_eclass
  mkeclass_axi4lite soc_eclass(.resetpc(64'd4096),
			       .CLK(CLK),
			       .RST_N(RST_N),
			       .master_d_m_arready_arready(soc_eclass_master_d_m_arready_arready),
			       .master_d_m_awready_awready(soc_eclass_master_d_m_awready_awready),
			       .master_d_m_bvalid_bresp(soc_eclass_master_d_m_bvalid_bresp),
			       .master_d_m_bvalid_bvalid(soc_eclass_master_d_m_bvalid_bvalid),
			       .master_d_m_rvalid_rdata(soc_eclass_master_d_m_rvalid_rdata),
			       .master_d_m_rvalid_rresp(soc_eclass_master_d_m_rvalid_rresp),
			       .master_d_m_rvalid_rvalid(soc_eclass_master_d_m_rvalid_rvalid),
			       .master_d_m_wready_wready(soc_eclass_master_d_m_wready_wready),
			       .master_i_m_arready_arready(soc_eclass_master_i_m_arready_arready),
			       .master_i_m_awready_awready(soc_eclass_master_i_m_awready_awready),
			       .master_i_m_bvalid_bresp(soc_eclass_master_i_m_bvalid_bresp),
			       .master_i_m_bvalid_bvalid(soc_eclass_master_i_m_bvalid_bvalid),
			       .master_i_m_rvalid_rdata(soc_eclass_master_i_m_rvalid_rdata),
			       .master_i_m_rvalid_rresp(soc_eclass_master_i_m_rvalid_rresp),
			       .master_i_m_rvalid_rvalid(soc_eclass_master_i_m_rvalid_rvalid),
			       .master_i_m_wready_wready(soc_eclass_master_i_m_wready_wready),
			       .sb_clint_msip_put(soc_eclass_sb_clint_msip_put),
			       .sb_clint_mtime_put(soc_eclass_sb_clint_mtime_put),
			       .sb_clint_mtip_put(soc_eclass_sb_clint_mtip_put),
			       .sb_ext_interrupt_put(soc_eclass_sb_ext_interrupt_put),
			       .EN_sb_clint_msip_put(soc_eclass_EN_sb_clint_msip_put),
			       .EN_sb_clint_mtip_put(soc_eclass_EN_sb_clint_mtip_put),
			       .EN_sb_clint_mtime_put(soc_eclass_EN_sb_clint_mtime_put),
			       .EN_sb_ext_interrupt_put(soc_eclass_EN_sb_ext_interrupt_put),
			       .EN_io_dump_get(soc_eclass_EN_io_dump_get),
			       .master_d_awvalid(soc_eclass_master_d_awvalid),
			       .master_d_awaddr(soc_eclass_master_d_awaddr),
			       .master_d_awprot(soc_eclass_master_d_awprot),
			       .master_d_awsize(soc_eclass_master_d_awsize),
			       .master_d_wvalid(soc_eclass_master_d_wvalid),
			       .master_d_wdata(soc_eclass_master_d_wdata),
			       .master_d_wstrb(soc_eclass_master_d_wstrb),
			       .master_d_bready(soc_eclass_master_d_bready),
			       .master_d_arvalid(soc_eclass_master_d_arvalid),
			       .master_d_araddr(soc_eclass_master_d_araddr),
			       .master_d_arprot(soc_eclass_master_d_arprot),
			       .master_d_arsize(soc_eclass_master_d_arsize),
			       .master_d_rready(soc_eclass_master_d_rready),
			       .master_i_awvalid(soc_eclass_master_i_awvalid),
			       .master_i_awaddr(soc_eclass_master_i_awaddr),
			       .master_i_awprot(soc_eclass_master_i_awprot),
			       .master_i_awsize(soc_eclass_master_i_awsize),
			       .master_i_wvalid(soc_eclass_master_i_wvalid),
			       .master_i_wdata(soc_eclass_master_i_wdata),
			       .master_i_wstrb(soc_eclass_master_i_wstrb),
			       .master_i_bready(soc_eclass_master_i_bready),
			       .master_i_arvalid(soc_eclass_master_i_arvalid),
			       .master_i_araddr(soc_eclass_master_i_araddr),
			       .master_i_arprot(soc_eclass_master_i_arprot),
			       .master_i_arsize(soc_eclass_master_i_arsize),
			       .master_i_rready(soc_eclass_master_i_rready),
			       .RDY_sb_clint_msip_put(),
			       .RDY_sb_clint_mtip_put(),
			       .RDY_sb_clint_mtime_put(),
			       .RDY_sb_ext_interrupt_put(),
			       .io_dump_get(),
			       .RDY_io_dump_get());

  // submodule soc_err_slave_s_xactor_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_err_slave_s_xactor_f_rd_addr(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(soc_err_slave_s_xactor_f_rd_addr_D_IN),
							    .ENQ(soc_err_slave_s_xactor_f_rd_addr_ENQ),
							    .DEQ(soc_err_slave_s_xactor_f_rd_addr_DEQ),
							    .CLR(soc_err_slave_s_xactor_f_rd_addr_CLR),
							    .D_OUT(),
							    .FULL_N(soc_err_slave_s_xactor_f_rd_addr_FULL_N),
							    .EMPTY_N(soc_err_slave_s_xactor_f_rd_addr_EMPTY_N));

  // submodule soc_err_slave_s_xactor_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_err_slave_s_xactor_f_rd_data(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(soc_err_slave_s_xactor_f_rd_data_D_IN),
							    .ENQ(soc_err_slave_s_xactor_f_rd_data_ENQ),
							    .DEQ(soc_err_slave_s_xactor_f_rd_data_DEQ),
							    .CLR(soc_err_slave_s_xactor_f_rd_data_CLR),
							    .D_OUT(soc_err_slave_s_xactor_f_rd_data_D_OUT),
							    .FULL_N(soc_err_slave_s_xactor_f_rd_data_FULL_N),
							    .EMPTY_N(soc_err_slave_s_xactor_f_rd_data_EMPTY_N));

  // submodule soc_err_slave_s_xactor_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_err_slave_s_xactor_f_wr_addr(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(soc_err_slave_s_xactor_f_wr_addr_D_IN),
							    .ENQ(soc_err_slave_s_xactor_f_wr_addr_ENQ),
							    .DEQ(soc_err_slave_s_xactor_f_wr_addr_DEQ),
							    .CLR(soc_err_slave_s_xactor_f_wr_addr_CLR),
							    .D_OUT(),
							    .FULL_N(soc_err_slave_s_xactor_f_wr_addr_FULL_N),
							    .EMPTY_N(soc_err_slave_s_xactor_f_wr_addr_EMPTY_N));

  // submodule soc_err_slave_s_xactor_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_err_slave_s_xactor_f_wr_data(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(soc_err_slave_s_xactor_f_wr_data_D_IN),
							    .ENQ(soc_err_slave_s_xactor_f_wr_data_ENQ),
							    .DEQ(soc_err_slave_s_xactor_f_wr_data_DEQ),
							    .CLR(soc_err_slave_s_xactor_f_wr_data_CLR),
							    .D_OUT(),
							    .FULL_N(soc_err_slave_s_xactor_f_wr_data_FULL_N),
							    .EMPTY_N(soc_err_slave_s_xactor_f_wr_data_EMPTY_N));

  // submodule soc_err_slave_s_xactor_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_err_slave_s_xactor_f_wr_resp(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(soc_err_slave_s_xactor_f_wr_resp_D_IN),
							    .ENQ(soc_err_slave_s_xactor_f_wr_resp_ENQ),
							    .DEQ(soc_err_slave_s_xactor_f_wr_resp_DEQ),
							    .CLR(soc_err_slave_s_xactor_f_wr_resp_CLR),
							    .D_OUT(soc_err_slave_s_xactor_f_wr_resp_D_OUT),
							    .FULL_N(soc_err_slave_s_xactor_f_wr_resp_FULL_N),
							    .EMPTY_N(soc_err_slave_s_xactor_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_v_f_rd_err_user_0
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_rd_err_user_0(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_rd_err_user_0_ENQ),
							 .DEQ(soc_fabric_v_f_rd_err_user_0_DEQ),
							 .CLR(soc_fabric_v_f_rd_err_user_0_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_rd_err_user_1
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_rd_err_user_1(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_rd_err_user_1_ENQ),
							 .DEQ(soc_fabric_v_f_rd_err_user_1_DEQ),
							 .CLR(soc_fabric_v_f_rd_err_user_1_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_rd_err_user_2
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_rd_err_user_2(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_rd_err_user_2_ENQ),
							 .DEQ(soc_fabric_v_f_rd_err_user_2_DEQ),
							 .CLR(soc_fabric_v_f_rd_err_user_2_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_rd_mis_0
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_0(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_0_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_0_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_0_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_0_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_0_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_0_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_0_EMPTY_N));

  // submodule soc_fabric_v_f_rd_mis_1
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_1(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_1_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_1_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_1_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_1_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_1_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_1_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_1_EMPTY_N));

  // submodule soc_fabric_v_f_rd_mis_2
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_2(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_2_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_2_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_2_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_2_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_2_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_2_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_2_EMPTY_N));

  // submodule soc_fabric_v_f_rd_mis_3
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_3(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_3_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_3_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_3_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_3_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_3_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_3_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_3_EMPTY_N));

  // submodule soc_fabric_v_f_rd_mis_4
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_4(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_4_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_4_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_4_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_4_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_4_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_4_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_4_EMPTY_N));

  // submodule soc_fabric_v_f_rd_mis_5
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_rd_mis_5(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_mis_5_D_IN),
								  .ENQ(soc_fabric_v_f_rd_mis_5_ENQ),
								  .DEQ(soc_fabric_v_f_rd_mis_5_DEQ),
								  .CLR(soc_fabric_v_f_rd_mis_5_CLR),
								  .D_OUT(soc_fabric_v_f_rd_mis_5_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_mis_5_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_mis_5_EMPTY_N));

  // submodule soc_fabric_v_f_rd_sjs_0
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_rd_sjs_0(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_sjs_0_D_IN),
								  .ENQ(soc_fabric_v_f_rd_sjs_0_ENQ),
								  .DEQ(soc_fabric_v_f_rd_sjs_0_DEQ),
								  .CLR(soc_fabric_v_f_rd_sjs_0_CLR),
								  .D_OUT(soc_fabric_v_f_rd_sjs_0_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_sjs_0_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_sjs_0_EMPTY_N));

  // submodule soc_fabric_v_f_rd_sjs_1
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_rd_sjs_1(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_sjs_1_D_IN),
								  .ENQ(soc_fabric_v_f_rd_sjs_1_ENQ),
								  .DEQ(soc_fabric_v_f_rd_sjs_1_DEQ),
								  .CLR(soc_fabric_v_f_rd_sjs_1_CLR),
								  .D_OUT(soc_fabric_v_f_rd_sjs_1_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_sjs_1_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_sjs_1_EMPTY_N));

  // submodule soc_fabric_v_f_rd_sjs_2
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_rd_sjs_2(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_rd_sjs_2_D_IN),
								  .ENQ(soc_fabric_v_f_rd_sjs_2_ENQ),
								  .DEQ(soc_fabric_v_f_rd_sjs_2_DEQ),
								  .CLR(soc_fabric_v_f_rd_sjs_2_CLR),
								  .D_OUT(soc_fabric_v_f_rd_sjs_2_D_OUT),
								  .FULL_N(soc_fabric_v_f_rd_sjs_2_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_rd_sjs_2_EMPTY_N));

  // submodule soc_fabric_v_f_wr_err_user_0
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_wr_err_user_0(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_wr_err_user_0_ENQ),
							 .DEQ(soc_fabric_v_f_wr_err_user_0_DEQ),
							 .CLR(soc_fabric_v_f_wr_err_user_0_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_wr_err_user_1
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_wr_err_user_1(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_wr_err_user_1_ENQ),
							 .DEQ(soc_fabric_v_f_wr_err_user_1_DEQ),
							 .CLR(soc_fabric_v_f_wr_err_user_1_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_wr_err_user_2
  FIFO20 #(.guarded(32'd1)) soc_fabric_v_f_wr_err_user_2(.RST(RST_N),
							 .CLK(CLK),
							 .ENQ(soc_fabric_v_f_wr_err_user_2_ENQ),
							 .DEQ(soc_fabric_v_f_wr_err_user_2_DEQ),
							 .CLR(soc_fabric_v_f_wr_err_user_2_CLR),
							 .FULL_N(),
							 .EMPTY_N());

  // submodule soc_fabric_v_f_wr_mis_0
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_0(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_0_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_0_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_0_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_0_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_0_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_0_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_0_EMPTY_N));

  // submodule soc_fabric_v_f_wr_mis_1
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_1(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_1_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_1_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_1_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_1_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_1_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_1_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_1_EMPTY_N));

  // submodule soc_fabric_v_f_wr_mis_2
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_2(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_2_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_2_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_2_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_2_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_2_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_2_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_2_EMPTY_N));

  // submodule soc_fabric_v_f_wr_mis_3
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_3(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_3_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_3_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_3_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_3_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_3_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_3_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_3_EMPTY_N));

  // submodule soc_fabric_v_f_wr_mis_4
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_4(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_4_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_4_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_4_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_4_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_4_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_4_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_4_EMPTY_N));

  // submodule soc_fabric_v_f_wr_mis_5
  FIFO2 #(.width(32'd2), .guarded(32'd1)) soc_fabric_v_f_wr_mis_5(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_mis_5_D_IN),
								  .ENQ(soc_fabric_v_f_wr_mis_5_ENQ),
								  .DEQ(soc_fabric_v_f_wr_mis_5_DEQ),
								  .CLR(soc_fabric_v_f_wr_mis_5_CLR),
								  .D_OUT(soc_fabric_v_f_wr_mis_5_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_mis_5_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_mis_5_EMPTY_N));

  // submodule soc_fabric_v_f_wr_sjs_0
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_wr_sjs_0(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_sjs_0_D_IN),
								  .ENQ(soc_fabric_v_f_wr_sjs_0_ENQ),
								  .DEQ(soc_fabric_v_f_wr_sjs_0_DEQ),
								  .CLR(soc_fabric_v_f_wr_sjs_0_CLR),
								  .D_OUT(soc_fabric_v_f_wr_sjs_0_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_sjs_0_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_sjs_0_EMPTY_N));

  // submodule soc_fabric_v_f_wr_sjs_1
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_wr_sjs_1(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_sjs_1_D_IN),
								  .ENQ(soc_fabric_v_f_wr_sjs_1_ENQ),
								  .DEQ(soc_fabric_v_f_wr_sjs_1_DEQ),
								  .CLR(soc_fabric_v_f_wr_sjs_1_CLR),
								  .D_OUT(soc_fabric_v_f_wr_sjs_1_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_sjs_1_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_sjs_1_EMPTY_N));

  // submodule soc_fabric_v_f_wr_sjs_2
  FIFO2 #(.width(32'd3), .guarded(32'd1)) soc_fabric_v_f_wr_sjs_2(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(soc_fabric_v_f_wr_sjs_2_D_IN),
								  .ENQ(soc_fabric_v_f_wr_sjs_2_ENQ),
								  .DEQ(soc_fabric_v_f_wr_sjs_2_DEQ),
								  .CLR(soc_fabric_v_f_wr_sjs_2_CLR),
								  .D_OUT(soc_fabric_v_f_wr_sjs_2_D_OUT),
								  .FULL_N(soc_fabric_v_f_wr_sjs_2_FULL_N),
								  .EMPTY_N(soc_fabric_v_f_wr_sjs_2_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_0_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_0_f_rd_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_0_f_rd_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_0_f_rd_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_0_f_rd_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_0_f_rd_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_0_f_rd_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_0_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_0_f_rd_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_0_f_rd_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_0_f_rd_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_0_f_rd_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_0_f_rd_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_0_f_rd_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_0_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_0_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_0_f_wr_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_0_f_wr_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_0_f_wr_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_0_f_wr_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_0_f_wr_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_0_f_wr_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_0_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_0_f_wr_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_0_f_wr_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_0_f_wr_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_0_f_wr_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_0_f_wr_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_0_f_wr_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_0_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_0_f_wr_resp(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_0_f_wr_resp_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_0_f_wr_resp_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_0_f_wr_resp_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_0_f_wr_resp_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_0_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_1_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_1_f_rd_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_1_f_rd_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_1_f_rd_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_1_f_rd_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_1_f_rd_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_1_f_rd_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_1_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_1_f_rd_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_1_f_rd_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_1_f_rd_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_1_f_rd_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_1_f_rd_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_1_f_rd_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_1_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_1_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_1_f_wr_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_1_f_wr_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_1_f_wr_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_1_f_wr_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_1_f_wr_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_1_f_wr_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_1_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_1_f_wr_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_1_f_wr_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_1_f_wr_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_1_f_wr_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_1_f_wr_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_1_f_wr_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_1_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_1_f_wr_resp(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_1_f_wr_resp_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_1_f_wr_resp_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_1_f_wr_resp_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_1_f_wr_resp_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_1_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_2_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_2_f_rd_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_2_f_rd_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_2_f_rd_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_2_f_rd_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_2_f_rd_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_2_f_rd_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_2_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_2_f_rd_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_2_f_rd_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_2_f_rd_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_2_f_rd_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_2_f_rd_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_2_f_rd_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_2_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_2_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_2_f_wr_addr(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_2_f_wr_addr_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_2_f_wr_addr_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_2_f_wr_addr_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_2_f_wr_addr_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_2_f_wr_addr_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_2_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_2_f_wr_data(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_2_f_wr_data_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_2_f_wr_data_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_2_f_wr_data_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_2_f_wr_data_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_2_f_wr_data_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_from_masters_2_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_from_masters_2_f_wr_resp(.RST(RST_N),
								       .CLK(CLK),
								       .D_IN(soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN),
								       .ENQ(soc_fabric_xactors_from_masters_2_f_wr_resp_ENQ),
								       .DEQ(soc_fabric_xactors_from_masters_2_f_wr_resp_DEQ),
								       .CLR(soc_fabric_xactors_from_masters_2_f_wr_resp_CLR),
								       .D_OUT(soc_fabric_xactors_from_masters_2_f_wr_resp_D_OUT),
								       .FULL_N(soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N),
								       .EMPTY_N(soc_fabric_xactors_from_masters_2_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_0_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_0_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_0_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_0_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_0_f_rd_addr_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_0_f_rd_addr_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_0_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_0_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_0_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_0_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_0_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_0_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT),
								    .FULL_N(),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_0_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_0_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_0_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_0_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_0_f_wr_addr_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_0_f_wr_addr_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_0_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_0_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_0_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_0_f_wr_data_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_0_f_wr_data_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_0_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_0_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_0_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_0_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_0_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT),
								    .FULL_N(),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_0_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_1_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_1_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_1_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_1_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_1_f_rd_addr_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_1_f_rd_addr_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_1_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_1_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_1_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_1_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_1_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_1_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT),
								    .FULL_N(),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_1_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_1_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_1_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_1_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_1_f_wr_addr_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_1_f_wr_addr_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_1_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_1_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_1_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_1_f_wr_data_CLR),
								    .D_OUT(),
								    .FULL_N(soc_fabric_xactors_to_slaves_1_f_wr_data_FULL_N),
								    .EMPTY_N());

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_1_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_1_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_1_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_1_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_1_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT),
								    .FULL_N(),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_1_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_2_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_2_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_2_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_2_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_2_f_rd_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_2_f_rd_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_2_f_rd_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_2_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_2_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_2_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_2_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_2_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_2_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_2_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_2_f_rd_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_2_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_2_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_2_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_2_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_2_f_wr_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_2_f_wr_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_2_f_wr_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_2_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_2_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_2_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_2_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_2_f_wr_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_2_f_wr_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_2_f_wr_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_2_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_2_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_2_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_2_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_2_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_2_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_2_f_wr_resp_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_2_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_3_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_3_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_3_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_3_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_3_f_rd_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_3_f_rd_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_3_f_rd_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_3_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_3_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_3_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_3_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_3_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_3_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_3_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_3_f_rd_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_3_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_3_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_3_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_3_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_3_f_wr_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_3_f_wr_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_3_f_wr_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_3_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_3_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_3_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_3_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_3_f_wr_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_3_f_wr_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_3_f_wr_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_3_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_3_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_3_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_3_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_3_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_3_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_3_f_wr_resp_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_3_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_4_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_4_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_4_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_4_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_4_f_rd_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_4_f_rd_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_4_f_rd_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_4_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_4_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_4_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_4_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_4_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_4_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_4_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_4_f_rd_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_4_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_4_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_4_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_4_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_4_f_wr_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_4_f_wr_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_4_f_wr_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_4_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_4_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_4_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_4_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_4_f_wr_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_4_f_wr_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_4_f_wr_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_4_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_4_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_4_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_4_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_4_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_4_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_4_f_wr_resp_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_4_f_wr_resp_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_5_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_5_f_rd_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_5_f_rd_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_5_f_rd_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_5_f_rd_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_5_f_rd_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_5_f_rd_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_5_f_rd_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_5_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_5_f_rd_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_5_f_rd_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_5_f_rd_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_5_f_rd_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_5_f_rd_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_5_f_rd_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_5_f_rd_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_5_f_wr_addr(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_5_f_wr_addr_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_5_f_wr_addr_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_5_f_wr_addr_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_5_f_wr_addr_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_5_f_wr_addr_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_5_f_wr_addr_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_5_f_wr_data(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_5_f_wr_data_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_5_f_wr_data_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_5_f_wr_data_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_5_f_wr_data_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_5_f_wr_data_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_5_f_wr_data_EMPTY_N));

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_fabric_xactors_to_slaves_5_f_wr_resp(.RST(RST_N),
								    .CLK(CLK),
								    .D_IN(soc_fabric_xactors_to_slaves_5_f_wr_resp_D_IN),
								    .ENQ(soc_fabric_xactors_to_slaves_5_f_wr_resp_ENQ),
								    .DEQ(soc_fabric_xactors_to_slaves_5_f_wr_resp_DEQ),
								    .CLR(soc_fabric_xactors_to_slaves_5_f_wr_resp_CLR),
								    .D_OUT(soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT),
								    .FULL_N(soc_fabric_xactors_to_slaves_5_f_wr_resp_FULL_N),
								    .EMPTY_N(soc_fabric_xactors_to_slaves_5_f_wr_resp_EMPTY_N));

  // submodule soc_signature
  mksign_dump_axi4lite soc_signature(.CLK(CLK),
				     .RST_N(RST_N),
				     .master_m_arready_arready(soc_signature_master_m_arready_arready),
				     .master_m_awready_awready(soc_signature_master_m_awready_awready),
				     .master_m_bvalid_bresp(soc_signature_master_m_bvalid_bresp),
				     .master_m_bvalid_bvalid(soc_signature_master_m_bvalid_bvalid),
				     .master_m_rvalid_rdata(soc_signature_master_m_rvalid_rdata),
				     .master_m_rvalid_rresp(soc_signature_master_m_rvalid_rresp),
				     .master_m_rvalid_rvalid(soc_signature_master_m_rvalid_rvalid),
				     .master_m_wready_wready(soc_signature_master_m_wready_wready),
				     .slave_m_arvalid_araddr(soc_signature_slave_m_arvalid_araddr),
				     .slave_m_arvalid_arprot(soc_signature_slave_m_arvalid_arprot),
				     .slave_m_arvalid_arsize(soc_signature_slave_m_arvalid_arsize),
				     .slave_m_arvalid_arvalid(soc_signature_slave_m_arvalid_arvalid),
				     .slave_m_awvalid_awaddr(soc_signature_slave_m_awvalid_awaddr),
				     .slave_m_awvalid_awprot(soc_signature_slave_m_awvalid_awprot),
				     .slave_m_awvalid_awsize(soc_signature_slave_m_awvalid_awsize),
				     .slave_m_awvalid_awvalid(soc_signature_slave_m_awvalid_awvalid),
				     .slave_m_bready_bready(soc_signature_slave_m_bready_bready),
				     .slave_m_rready_rready(soc_signature_slave_m_rready_rready),
				     .slave_m_wvalid_wdata(soc_signature_slave_m_wvalid_wdata),
				     .slave_m_wvalid_wstrb(soc_signature_slave_m_wvalid_wstrb),
				     .slave_m_wvalid_wvalid(soc_signature_slave_m_wvalid_wvalid),
				     .master_awvalid(soc_signature_master_awvalid),
				     .master_awaddr(soc_signature_master_awaddr),
				     .master_awprot(soc_signature_master_awprot),
				     .master_awsize(soc_signature_master_awsize),
				     .master_wvalid(soc_signature_master_wvalid),
				     .master_wdata(soc_signature_master_wdata),
				     .master_wstrb(soc_signature_master_wstrb),
				     .master_bready(soc_signature_master_bready),
				     .master_arvalid(soc_signature_master_arvalid),
				     .master_araddr(soc_signature_master_araddr),
				     .master_arprot(soc_signature_master_arprot),
				     .master_arsize(soc_signature_master_arsize),
				     .master_rready(soc_signature_master_rready),
				     .slave_awready(soc_signature_slave_awready),
				     .slave_wready(soc_signature_slave_wready),
				     .slave_bvalid(soc_signature_slave_bvalid),
				     .slave_bresp(soc_signature_slave_bresp),
				     .slave_arready(soc_signature_slave_arready),
				     .slave_rvalid(soc_signature_slave_rvalid),
				     .slave_rresp(soc_signature_slave_rresp),
				     .slave_rdata(soc_signature_slave_rdata),
				     .mv_end_simulation(),
				     .RDY_mv_end_simulation());

  // submodule soc_uart_s_xactor_f_rd_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_uart_s_xactor_f_rd_addr(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(soc_uart_s_xactor_f_rd_addr_D_IN),
						       .ENQ(soc_uart_s_xactor_f_rd_addr_ENQ),
						       .DEQ(soc_uart_s_xactor_f_rd_addr_DEQ),
						       .CLR(soc_uart_s_xactor_f_rd_addr_CLR),
						       .D_OUT(soc_uart_s_xactor_f_rd_addr_D_OUT),
						       .FULL_N(soc_uart_s_xactor_f_rd_addr_FULL_N),
						       .EMPTY_N(soc_uart_s_xactor_f_rd_addr_EMPTY_N));

  // submodule soc_uart_s_xactor_f_rd_data
  FIFO2 #(.width(32'd66),
	  .guarded(32'd1)) soc_uart_s_xactor_f_rd_data(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(soc_uart_s_xactor_f_rd_data_D_IN),
						       .ENQ(soc_uart_s_xactor_f_rd_data_ENQ),
						       .DEQ(soc_uart_s_xactor_f_rd_data_DEQ),
						       .CLR(soc_uart_s_xactor_f_rd_data_CLR),
						       .D_OUT(soc_uart_s_xactor_f_rd_data_D_OUT),
						       .FULL_N(soc_uart_s_xactor_f_rd_data_FULL_N),
						       .EMPTY_N(soc_uart_s_xactor_f_rd_data_EMPTY_N));

  // submodule soc_uart_s_xactor_f_wr_addr
  FIFO2 #(.width(32'd37),
	  .guarded(32'd1)) soc_uart_s_xactor_f_wr_addr(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(soc_uart_s_xactor_f_wr_addr_D_IN),
						       .ENQ(soc_uart_s_xactor_f_wr_addr_ENQ),
						       .DEQ(soc_uart_s_xactor_f_wr_addr_DEQ),
						       .CLR(soc_uart_s_xactor_f_wr_addr_CLR),
						       .D_OUT(soc_uart_s_xactor_f_wr_addr_D_OUT),
						       .FULL_N(soc_uart_s_xactor_f_wr_addr_FULL_N),
						       .EMPTY_N(soc_uart_s_xactor_f_wr_addr_EMPTY_N));

  // submodule soc_uart_s_xactor_f_wr_data
  FIFO2 #(.width(32'd72),
	  .guarded(32'd1)) soc_uart_s_xactor_f_wr_data(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(soc_uart_s_xactor_f_wr_data_D_IN),
						       .ENQ(soc_uart_s_xactor_f_wr_data_ENQ),
						       .DEQ(soc_uart_s_xactor_f_wr_data_DEQ),
						       .CLR(soc_uart_s_xactor_f_wr_data_CLR),
						       .D_OUT(soc_uart_s_xactor_f_wr_data_D_OUT),
						       .FULL_N(soc_uart_s_xactor_f_wr_data_FULL_N),
						       .EMPTY_N(soc_uart_s_xactor_f_wr_data_EMPTY_N));

  // submodule soc_uart_s_xactor_f_wr_resp
  FIFO2 #(.width(32'd2),
	  .guarded(32'd1)) soc_uart_s_xactor_f_wr_resp(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(soc_uart_s_xactor_f_wr_resp_D_IN),
						       .ENQ(soc_uart_s_xactor_f_wr_resp_ENQ),
						       .DEQ(soc_uart_s_xactor_f_wr_resp_DEQ),
						       .CLR(soc_uart_s_xactor_f_wr_resp_CLR),
						       .D_OUT(soc_uart_s_xactor_f_wr_resp_D_OUT),
						       .FULL_N(soc_uart_s_xactor_f_wr_resp_FULL_N),
						       .EMPTY_N(soc_uart_s_xactor_f_wr_resp_EMPTY_N));

  // submodule soc_uart_user_ifc_uart_baudGen_rBaudCounter
  Counter #(.width(32'd16),
	    .init(16'd0)) soc_uart_user_ifc_uart_baudGen_rBaudCounter(.CLK(CLK),
								      .RST(RST_N),
								      .DATA_A(soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_A),
								      .DATA_B(soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_B),
								      .DATA_C(soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_C),
								      .DATA_F(soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_F),
								      .ADDA(soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDA),
								      .ADDB(soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDB),
								      .SETC(soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETC),
								      .SETF(soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETF),
								      .Q_OUT(soc_uart_user_ifc_uart_baudGen_rBaudCounter_Q_OUT));

  // submodule soc_uart_user_ifc_uart_baudGen_rBaudTickCounter
  Counter #(.width(32'd3),
	    .init(3'd0)) soc_uart_user_ifc_uart_baudGen_rBaudTickCounter(.CLK(CLK),
									 .RST(RST_N),
									 .DATA_A(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_A),
									 .DATA_B(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_B),
									 .DATA_C(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_C),
									 .DATA_F(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_F),
									 .ADDA(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDA),
									 .ADDB(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDB),
									 .SETC(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETC),
									 .SETF(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETF),
									 .Q_OUT(soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_Q_OUT));

  // submodule soc_uart_user_ifc_uart_fifoRecv
  SizedFIFO #(.p1width(32'd8),
	      .p2depth(32'd16),
	      .p3cntr_width(32'd4),
	      .guarded(32'd1)) soc_uart_user_ifc_uart_fifoRecv(.RST(RST_N),
							       .CLK(CLK),
							       .D_IN(soc_uart_user_ifc_uart_fifoRecv_D_IN),
							       .ENQ(soc_uart_user_ifc_uart_fifoRecv_ENQ),
							       .DEQ(soc_uart_user_ifc_uart_fifoRecv_DEQ),
							       .CLR(soc_uart_user_ifc_uart_fifoRecv_CLR),
							       .D_OUT(soc_uart_user_ifc_uart_fifoRecv_D_OUT),
							       .FULL_N(soc_uart_user_ifc_uart_fifoRecv_FULL_N),
							       .EMPTY_N(soc_uart_user_ifc_uart_fifoRecv_EMPTY_N));

  // submodule soc_uart_user_ifc_uart_fifoXmit
  SizedFIFO #(.p1width(32'd8),
	      .p2depth(32'd16),
	      .p3cntr_width(32'd4),
	      .guarded(32'd1)) soc_uart_user_ifc_uart_fifoXmit(.RST(RST_N),
							       .CLK(CLK),
							       .D_IN(soc_uart_user_ifc_uart_fifoXmit_D_IN),
							       .ENQ(soc_uart_user_ifc_uart_fifoXmit_ENQ),
							       .DEQ(soc_uart_user_ifc_uart_fifoXmit_DEQ),
							       .CLR(soc_uart_user_ifc_uart_fifoXmit_CLR),
							       .D_OUT(soc_uart_user_ifc_uart_fifoXmit_D_OUT),
							       .FULL_N(soc_uart_user_ifc_uart_fifoXmit_FULL_N),
							       .EMPTY_N(soc_uart_user_ifc_uart_fifoXmit_EMPTY_N));

  // rule RL_soc_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_FULL_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_1
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16) &&
	     !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_2
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d51 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_3
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_FULL_N &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16) &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d68 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_4
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d88 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_5
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d103 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_6
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 =
	     soc_fabric_xactors_to_slaves_0_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_7
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 =
	     soc_fabric_xactors_to_slaves_1_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117) &&
	     !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_8
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 =
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d142 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_9
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 =
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117) &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d154 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_10
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d169 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_11
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 =
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d179 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_12
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 =
	     soc_fabric_xactors_to_slaves_0_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_13
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 =
	     soc_fabric_xactors_to_slaves_1_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193) &&
	     !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_14
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 =
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d218 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_15
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 =
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193) &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d230 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_16
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d245 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_wr_xaction_master_to_slave_17
  assign CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 =
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_FULL_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_data_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d255 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 &&
	     !WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_FULL_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_1
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_1_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268) &&
	     !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_2
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d296 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_3
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_FULL_N &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268) &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d310 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_4
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d327 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_5
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_FULL_N &&
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d339 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_6
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 =
	     soc_fabric_xactors_to_slaves_0_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_7
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 =
	     soc_fabric_xactors_to_slaves_1_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350) &&
	     !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_8
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 =
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d372 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_9
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 =
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350) &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d383 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_10
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d397 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_11
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 =
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_FULL_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d406 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_12
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 =
	     soc_fabric_xactors_to_slaves_0_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_13
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 =
	     soc_fabric_xactors_to_slaves_1_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417) &&
	     !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_14
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 =
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d439 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_15
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 =
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417) &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d450 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_16
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d464 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ;

  // rule RL_soc_fabric_rl_rd_xaction_master_to_slave_17
  assign CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 =
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_FULL_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d473 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 &&
	     !WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master =
	     soc_fabric_v_f_wr_mis_0_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_resp_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_1
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 =
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_mis_1_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_2
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 =
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_mis_2_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_3
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 =
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_mis_3_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_4
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 =
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_mis_4_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_5
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 =
	     soc_fabric_v_f_wr_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_mis_5_D_OUT == 2'd0 &&
	     soc_fabric_v_f_wr_sjs_0_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_6
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 =
	     soc_fabric_v_f_wr_mis_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_7
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 =
	     soc_fabric_v_f_wr_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_8
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 =
	     soc_fabric_v_f_wr_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_9
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 =
	     soc_fabric_v_f_wr_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_10
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 =
	     soc_fabric_v_f_wr_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_11
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 =
	     soc_fabric_v_f_wr_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_D_OUT == 2'd1 &&
	     soc_fabric_v_f_wr_sjs_1_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_12
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 =
	     soc_fabric_v_f_wr_mis_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_0_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_13
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 =
	     soc_fabric_v_f_wr_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_1_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_14
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 =
	     soc_fabric_v_f_wr_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_2_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_15
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 =
	     soc_fabric_v_f_wr_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_3_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_16
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 =
	     soc_fabric_v_f_wr_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_4_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 ;

  // rule RL_soc_fabric_rl_wr_resp_slave_to_master_17
  assign CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 =
	     soc_fabric_v_f_wr_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_resp_EMPTY_N &&
	     soc_fabric_v_f_wr_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_FULL_N &&
	     soc_fabric_v_f_wr_mis_5_D_OUT == 2'd2 &&
	     soc_fabric_v_f_wr_sjs_2_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 =
	     CAN_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master =
	     soc_fabric_v_f_rd_mis_0_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_rd_data_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_1
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 =
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_mis_1_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_2
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 =
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_mis_2_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_3
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 =
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_mis_3_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_4
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 =
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_mis_4_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_5
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 =
	     soc_fabric_v_f_rd_sjs_0_EMPTY_N &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_mis_5_D_OUT == 2'd0 &&
	     soc_fabric_v_f_rd_sjs_0_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_6
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 =
	     soc_fabric_v_f_rd_mis_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_7
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 =
	     soc_fabric_v_f_rd_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_8
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 =
	     soc_fabric_v_f_rd_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_9
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 =
	     soc_fabric_v_f_rd_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_10
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 =
	     soc_fabric_v_f_rd_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_11
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 =
	     soc_fabric_v_f_rd_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_1_EMPTY_N &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_D_OUT == 2'd1 &&
	     soc_fabric_v_f_rd_sjs_1_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_12
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 =
	     soc_fabric_v_f_rd_mis_0_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_0_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_0_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd0 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_13
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 =
	     soc_fabric_v_f_rd_mis_1_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_1_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_1_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd1 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_14
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 =
	     soc_fabric_v_f_rd_mis_2_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_2_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd2 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_15
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 =
	     soc_fabric_v_f_rd_mis_3_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_3_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd3 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_16
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 =
	     soc_fabric_v_f_rd_mis_4_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_4_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_4_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd4 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 ;

  // rule RL_soc_fabric_rl_rd_resp_slave_to_master_17
  assign CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 =
	     soc_fabric_v_f_rd_mis_5_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_rd_data_EMPTY_N &&
	     soc_fabric_v_f_rd_sjs_2_EMPTY_N &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_FULL_N &&
	     soc_fabric_v_f_rd_mis_5_D_OUT == 2'd2 &&
	     soc_fabric_v_f_rd_sjs_2_D_OUT == 3'd5 ;
  assign WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 =
	     CAN_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 ;

  // rule RL_soc_uart_user_ifc_capture_status
  assign CAN_FIRE_RL_soc_uart_user_ifc_capture_status = 1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_capture_status = 1'd1 ;

  // rule RL_soc_uart_capture_read_request
  assign CAN_FIRE_RL_soc_uart_capture_read_request =
	     soc_uart_s_xactor_f_rd_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_rd_data_FULL_N ;
  assign WILL_FIRE_RL_soc_uart_capture_read_request =
	     CAN_FIRE_RL_soc_uart_capture_read_request ;

  // rule RL_soc_uart_user_ifc_uart_baudGen_baud_count_wire
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_count_wire = 1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_count_wire = 1'd1 ;

  // rule RL_soc_uart_user_ifc_uart_baud_generator_clock_enable
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_baud_generator_clock_enable =
	     1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_baud_generator_clock_enable =
	     1'd1 ;

  // rule RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit =
	     soc_uart_user_ifc_uart_rRecvState == 3'd0 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit ;

  // rule RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell =
	     soc_uart_user_ifc_uart_rRecvState == 3'd1 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell ;

  // rule RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample =
	     soc_uart_user_ifc_uart_rRecvState == 3'd2 &&
	     soc_uart_user_ifc_uart_rRecvCellCount == 4'hF &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample ;

  // rule RL_soc_uart_user_ifc_uart_receive_sample_pin
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // rule RL_soc_uart_user_ifc_uart_receive_parity_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit =
	     soc_uart_user_ifc_uart_rRecvState == 3'd4 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ;

  // rule RL_soc_uart_user_ifc_uart_receive_stop_first_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit =
	     soc_uart_user_ifc_uart_rRecvState == 3'd5 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit ;

  // rule RL_soc_uart_user_ifc_uart_receive_bit_counter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_counter = 1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_counter = 1'd1 ;

  // rule RL_soc_uart_user_ifc_uart_receive_stop_last_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit =
	     soc_uart_user_ifc_uart_rRecvState == 3'd6 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit ;

  // rule RL_soc_uart_user_ifc_uart_receive_bit_cell_time_counter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_cell_time_counter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_bit_cell_time_counter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // rule RL_soc_uart_user_ifc_uart_receive_buffer_shift
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift =
	     soc_uart_user_ifc_uart_rRecvState == 3'd3 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // rule RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command =
	     soc_uart_user_ifc_uart_rXmitState == 3'd0 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ;

  // rule RL_soc_uart_capture_write_request
  assign CAN_FIRE_RL_soc_uart_capture_write_request =
	     soc_uart_s_xactor_f_wr_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_data_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_resp_FULL_N ;
  assign WILL_FIRE_RL_soc_uart_capture_write_request =
	     CAN_FIRE_RL_soc_uart_capture_write_request ;

  // rule RL_soc_uart_user_ifc_uart_transmit_send_start_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit =
	     soc_uart_user_ifc_uart_rXmitState == 3'd1 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit ;

  // rule RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time =
	     soc_uart_user_ifc_uart_rXmitState == 3'd2 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time ;

  // rule RL_soc_uart_user_ifc_uart_transmit_bit_counter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_counter = 1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_counter = 1'd1 ;

  // rule RL_soc_uart_user_ifc_uart_transmit_shift_next_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit =
	     soc_uart_user_ifc_uart_rXmitState == 3'd3 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit ;

  // rule RL_soc_uart_user_ifc_uart_transmit_buffer_load
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load =
	     soc_uart_user_ifc_uart_fifoXmit_EMPTY_N &&
	     soc_uart_user_ifc_uart_pwXmitLoadBuffer_whas ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ;

  // rule RL_soc_uart_user_ifc_uart_transmit_buffer_shift
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift =
	     !soc_uart_user_ifc_uart_pwXmitLoadBuffer_whas &&
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // rule RL_soc_uart_user_ifc_uart_transmit_send_parity_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit =
	     soc_uart_user_ifc_uart_rXmitState == 3'd7 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit ;

  // rule RL_soc_uart_user_ifc_uart_transmit_send_stop_bit
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit =
	     soc_uart_user_ifc_uart_rXmitState == 3'd4 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit ;

  // rule RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 =
	     soc_uart_user_ifc_uart_rXmitState == 3'd5 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 ;

  // rule RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 =
	     soc_uart_user_ifc_uart_rXmitState == 3'd6 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 ;

  // rule RL_soc_uart_user_ifc_uart_transmit_bit_cell_time_counter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_cell_time_counter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_bit_cell_time_counter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // rule RL_soc_uart_user_ifc_uart_baudGen_baud_tick_count_wire
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_tick_count_wire =
	     1'd1 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_baud_tick_count_wire =
	     1'd1 ;

  // rule RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick =
	     soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_Q_OUT == 3'd0 &&
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_assert_2x_baud_tick ;

  // rule RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x =
	     !soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // rule RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit !=
	     soc_uart_user_ifc_uart_fifoRecv_r_deq_whas ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter ;

  // rule RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter
  assign CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter =
	     soc_uart_user_ifc_uart_fifoXmit_r_enq_whas !=
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ;
  assign WILL_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter ;

  // rule RL_soc_clint_axi_read_transaction
  assign CAN_FIRE_RL_soc_clint_axi_read_transaction =
	     soc_clint_s_xactor_f_rd_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_rd_data_FULL_N ;
  assign WILL_FIRE_RL_soc_clint_axi_read_transaction =
	     CAN_FIRE_RL_soc_clint_axi_read_transaction ;

  // rule RL_soc_err_slave_receive_read_request
  assign CAN_FIRE_RL_soc_err_slave_receive_read_request =
	     soc_err_slave_s_xactor_f_rd_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_rd_data_FULL_N ;
  assign WILL_FIRE_RL_soc_err_slave_receive_read_request =
	     CAN_FIRE_RL_soc_err_slave_receive_read_request ;

  // rule RL_soc_err_slave_receive_write_request
  assign CAN_FIRE_RL_soc_err_slave_receive_write_request =
	     soc_err_slave_s_xactor_f_wr_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_data_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_resp_FULL_N ;
  assign WILL_FIRE_RL_soc_err_slave_receive_write_request =
	     CAN_FIRE_RL_soc_err_slave_receive_write_request ;

  // rule RL_soc_1_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_1_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_1_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_1_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_1_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_1_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_1_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_1_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_1_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_1_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_1_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_1_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_1_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_1_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_1_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_2_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_2_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_2_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_2_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_2_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_2_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_2_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_2_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_2_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_2_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_2_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_2_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_2_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_2_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_2_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_3_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_3_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_3_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_3_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_3_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_3_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_3_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_3_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_3_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_3_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_3_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_3_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_3_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_3_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_3_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_4_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_4_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_4_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_4_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_4_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_4_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_4_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_4_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_4_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_4_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_4_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_4_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_4_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_4_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_4_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_5_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_5_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_5_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_5_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_5_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_5_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_5_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_5_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_5_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_5_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_5_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_5_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_5_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_5_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_5_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_6_rl_wr_addr_channel
  assign CAN_FIRE_RL_soc_6_rl_wr_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_6_rl_wr_addr_channel = 1'd1 ;

  // rule RL_soc_6_rl_wr_data_channel
  assign CAN_FIRE_RL_soc_6_rl_wr_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_6_rl_wr_data_channel = 1'd1 ;

  // rule RL_soc_6_rl_wr_response_channel
  assign CAN_FIRE_RL_soc_6_rl_wr_response_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_6_rl_wr_response_channel = 1'd1 ;

  // rule RL_soc_6_rl_rd_addr_channel
  assign CAN_FIRE_RL_soc_6_rl_rd_addr_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_6_rl_rd_addr_channel = 1'd1 ;

  // rule RL_soc_6_rl_rd_data_channel
  assign CAN_FIRE_RL_soc_6_rl_rd_data_channel = 1'd1 ;
  assign WILL_FIRE_RL_soc_6_rl_rd_data_channel = 1'd1 ;

  // rule RL_soc_7_mkConnectionGetPut
  assign CAN_FIRE_RL_soc_7_mkConnectionGetPut = 1'd1 ;
  assign WILL_FIRE_RL_soc_7_mkConnectionGetPut = 1'd1 ;

  // rule RL_soc_clint_axi_write_transaction
  assign CAN_FIRE_RL_soc_clint_axi_write_transaction =
	     soc_clint_s_xactor_f_wr_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_data_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_resp_FULL_N ;
  assign WILL_FIRE_RL_soc_clint_axi_write_transaction =
	     CAN_FIRE_RL_soc_clint_axi_write_transaction ;

  // rule RL_soc_8_mkConnectionGetPut
  assign CAN_FIRE_RL_soc_8_mkConnectionGetPut = 1'd1 ;
  assign WILL_FIRE_RL_soc_8_mkConnectionGetPut = 1'd1 ;

  // rule RL_soc_clint_clint_generate_time_interrupt
  assign CAN_FIRE_RL_soc_clint_clint_generate_time_interrupt =
	     !soc_clint_clint_wr_mtimecmp_written_whas ;
  assign WILL_FIRE_RL_soc_clint_clint_generate_time_interrupt =
	     CAN_FIRE_RL_soc_clint_clint_generate_time_interrupt &&
	     !WILL_FIRE_RL_soc_clint_axi_write_transaction ;

  // rule RL_soc_clint_clint_clear_interrupt
  assign CAN_FIRE_RL_soc_clint_clint_clear_interrupt =
	     soc_clint_clint_wr_mtimecmp_written_whas ;
  assign WILL_FIRE_RL_soc_clint_clint_clear_interrupt =
	     soc_clint_clint_wr_mtimecmp_written_whas ;

  // rule RL_soc_9_mkConnectionGetPut
  assign CAN_FIRE_RL_soc_9_mkConnectionGetPut = 1'd1 ;
  assign WILL_FIRE_RL_soc_9_mkConnectionGetPut = 1'd1 ;

  // rule RL_soc_clint_clint_increment_timer
  assign CAN_FIRE_RL_soc_clint_clint_increment_timer = 1'd1 ;
  assign WILL_FIRE_RL_soc_clint_clint_increment_timer = 1'd1 ;

  // inputs to muxes for submodule ports
  assign MUX_soc_uart_user_ifc_uart_rRecvState_write_1__SEL_6 =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin ;
  assign MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_1 =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time ;
  assign MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_2 =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit ;
  assign MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_3 =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ;
  assign MUX_soc_clint_clint_mtip_write_1__VAL_1 =
	     soc_clint_clint_rgmtime >= soc_clint_clint_rgmtimecmp ;
  assign MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_1 =
	     soc_uart_user_ifc_uart_rRecvData ? 3'd0 : 3'd1 ;
  assign MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_2 =
	     (soc_uart_user_ifc_uart_rRecvCellCount == 4'h4) ?
	       (soc_uart_user_ifc_uart_rRecvData ? 3'd0 : 3'd2) :
	       3'd1 ;
  always@(soc_uart_user_ifc_uart_rRecvBitCount)
  begin
    case (soc_uart_user_ifc_uart_rRecvBitCount)
      4'd8, 4'd9, 4'd10:
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_3 = 3'd6;
      default: MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_3 = 3'd3;
    endcase
  end
  assign MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_4 =
	     soc_uart_user_ifc_uart_rRecvData ? 3'd2 : 3'd0 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_1 =
	     soc_uart_user_ifc_uart_fifoXmit_EMPTY_N ? 3'd1 : 3'd0 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_2 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'hF) ? 3'd2 : 3'd1 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_3 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'hF) ?
	       ((soc_uart_user_ifc_uart_rXmitBitCount == 4'd7) ?
		  3'd4 :
		  3'd3) :
	       3'd2 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_4 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'hF) ? 3'd4 : 3'd7 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_5 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'hF) ? 3'd0 : 3'd4 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_6 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'h7) ? 3'd0 : 3'd5 ;
  assign MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_7 =
	     (soc_uart_user_ifc_uart_rXmitCellCount == 4'hF) ? 3'd0 : 3'd6 ;

  // inlined wires
  assign soc_uart_user_ifc_wr_status_wget =
	     { soc_uart_user_ifc_uart_fifoRecv_EMPTY_N,
	       soc_uart_user_ifc_uart_fifoRecv_FULL_N,
	       soc_uart_user_ifc_uart_fifoXmit_FULL_N,
	       !soc_uart_user_ifc_uart_fifoXmit_EMPTY_N &&
	       soc_uart_user_ifc_uart_rXmitState == 3'd0 } ;
  assign soc_clint_clint_wr_mtimecmp_written_whas =
	     WILL_FIRE_RL_soc_clint_axi_write_transaction &&
	     soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] >= 16'h4000 &&
	     soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] <= 16'd16391 ;
  assign soc_uart_user_ifc_uart_fifoRecv_r_deq_whas =
	     WILL_FIRE_RL_soc_uart_capture_read_request &&
	     soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'h8 &&
	     soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0 ;
  assign soc_uart_user_ifc_uart_pwRecvCellCountReset_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell &&
	     soc_uart_user_ifc_uart_rRecvCellCount == 4'h4 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit ;
  assign soc_uart_user_ifc_uart_pwRecvResetBitCount_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit &&
	     soc_uart_user_ifc_uart_rRecvData ;
  assign soc_uart_user_ifc_uart_pwRecvEnableBitCount_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin ;
  assign soc_uart_user_ifc_uart_fifoXmit_r_enq_whas =
	     WILL_FIRE_RL_soc_uart_capture_write_request &&
	     soc_uart_s_xactor_f_wr_addr_D_OUT[8:5] == 4'h4 &&
	     soc_uart_s_xactor_f_wr_addr_D_OUT[1:0] == 2'd0 ;
  assign soc_uart_user_ifc_uart_pwXmitCellCountReset_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command &&
	     soc_uart_user_ifc_uart_fifoXmit_EMPTY_N ||
	     _dor2soc_uart_user_ifc_uart_pwXmitCellCountReset_EN_wset &&
	     soc_uart_user_ifc_uart_rXmitCellCount == 4'hF ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 &&
	     soc_uart_user_ifc_uart_rXmitCellCount == 4'h7 ;
  assign soc_uart_user_ifc_uart_pwXmitEnableBitCount_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time &&
	     soc_uart_user_ifc_uart_rXmitCellCount == 4'hF &&
	     soc_uart_user_ifc_uart_rXmitBitCount != 4'd7 ;
  assign soc_uart_user_ifc_uart_pwXmitLoadBuffer_whas =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command &&
	     soc_uart_user_ifc_uart_fifoXmit_EMPTY_N ;

  // register soc_clint_clint_msip
  assign soc_clint_clint_msip_D_IN = data__h56748[0] ;
  assign soc_clint_clint_msip_EN =
	     WILL_FIRE_RL_soc_clint_axi_write_transaction &&
	     soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] == 16'h0 ;

  // register soc_clint_clint_mtip
  assign soc_clint_clint_mtip_D_IN =
	     WILL_FIRE_RL_soc_clint_clint_generate_time_interrupt &&
	     MUX_soc_clint_clint_mtip_write_1__VAL_1 ;
  assign soc_clint_clint_mtip_EN =
	     WILL_FIRE_RL_soc_clint_clint_generate_time_interrupt ||
	     soc_clint_clint_wr_mtimecmp_written_whas ;

  // register soc_clint_clint_rg_tick
  assign soc_clint_clint_rg_tick_D_IN = soc_clint_clint_rg_tick + 4'd1 ;
  assign soc_clint_clint_rg_tick_EN = 1'd1 ;

  // register soc_clint_clint_rgmtime
  assign soc_clint_clint_rgmtime_D_IN = soc_clint_clint_rgmtime + 64'd1 ;
  assign soc_clint_clint_rgmtime_EN = soc_clint_clint_rg_tick == 4'd0 ;

  // register soc_clint_clint_rgmtimecmp
  assign soc_clint_clint_rgmtimecmp_D_IN = x__h58828 | datamask__h56751 ;
  assign soc_clint_clint_rgmtimecmp_EN =
	     soc_clint_clint_wr_mtimecmp_written_whas ;

  // register soc_uart_user_ifc_baud_value
  assign soc_uart_user_ifc_baud_value_D_IN =
	     soc_uart_s_xactor_f_wr_data_D_OUT[23:8] ;
  assign soc_uart_user_ifc_baud_value_EN =
	     WILL_FIRE_RL_soc_uart_capture_write_request &&
	     soc_uart_s_xactor_f_wr_addr_D_OUT[8:5] == 4'h0 &&
	     soc_uart_s_xactor_f_wr_addr_D_OUT[1:0] == 2'd1 ;

  // register soc_uart_user_ifc_uart_fifoRecv_countReg
  assign soc_uart_user_ifc_uart_fifoRecv_countReg_D_IN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit ?
	       soc_uart_user_ifc_uart_fifoRecv_countReg + 5'd1 :
	       soc_uart_user_ifc_uart_fifoRecv_countReg - 5'd1 ;
  assign soc_uart_user_ifc_uart_fifoRecv_countReg_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoRecv__updateLevelCounter ;

  // register soc_uart_user_ifc_uart_fifoXmit_countReg
  assign soc_uart_user_ifc_uart_fifoXmit_countReg_D_IN =
	     soc_uart_user_ifc_uart_fifoXmit_r_enq_whas ?
	       soc_uart_user_ifc_uart_fifoXmit_countReg + 5'd1 :
	       soc_uart_user_ifc_uart_fifoXmit_countReg - 5'd1 ;
  assign soc_uart_user_ifc_uart_fifoXmit_countReg_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_fifoXmit__updateLevelCounter ;

  // register soc_uart_user_ifc_uart_rRecvBitCount
  assign soc_uart_user_ifc_uart_rRecvBitCount_D_IN =
	     soc_uart_user_ifc_uart_pwRecvResetBitCount_whas ?
	       4'd0 :
	       x__h35390 ;
  assign soc_uart_user_ifc_uart_rRecvBitCount_EN =
	     soc_uart_user_ifc_uart_pwRecvResetBitCount_whas ||
	     soc_uart_user_ifc_uart_pwRecvEnableBitCount_whas ;

  // register soc_uart_user_ifc_uart_rRecvCellCount
  assign soc_uart_user_ifc_uart_rRecvCellCount_D_IN =
	     soc_uart_user_ifc_uart_pwRecvCellCountReset_whas ?
	       4'd0 :
	       x__h33749 ;
  assign soc_uart_user_ifc_uart_rRecvCellCount_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // register soc_uart_user_ifc_uart_rRecvData
  assign soc_uart_user_ifc_uart_rRecvData_D_IN = 1'b0 ;
  assign soc_uart_user_ifc_uart_rRecvData_EN = 1'b0 ;

  // register soc_uart_user_ifc_uart_rRecvParity
  assign soc_uart_user_ifc_uart_rRecvParity_D_IN =
	     soc_uart_user_ifc_uart_rRecvData ;
  assign soc_uart_user_ifc_uart_rRecvParity_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ;

  // register soc_uart_user_ifc_uart_rRecvState
  always@(WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit or
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_1 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell or
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_2 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample or
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_3 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit or
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_4 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit or
	  MUX_soc_uart_user_ifc_uart_rRecvState_write_1__SEL_6)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit:
	  soc_uart_user_ifc_uart_rRecvState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_1;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell:
	  soc_uart_user_ifc_uart_rRecvState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_2;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample:
	  soc_uart_user_ifc_uart_rRecvState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_3;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit:
	  soc_uart_user_ifc_uart_rRecvState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rRecvState_write_1__VAL_4;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit:
	  soc_uart_user_ifc_uart_rRecvState_D_IN = 3'd0;
      MUX_soc_uart_user_ifc_uart_rRecvState_write_1__SEL_6:
	  soc_uart_user_ifc_uart_rRecvState_D_IN = 3'd2;
      default: soc_uart_user_ifc_uart_rRecvState_D_IN =
		   3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_uart_user_ifc_uart_rRecvState_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_for_start_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_find_center_of_bit_cell ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_wait_bit_cell_time_for_sample ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_first_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_receive_sample_pin ;

  // register soc_uart_user_ifc_uart_rXmitBitCount
  assign soc_uart_user_ifc_uart_rXmitBitCount_D_IN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ?
	       4'd0 :
	       x__h37208 ;
  assign soc_uart_user_ifc_uart_rXmitBitCount_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ||
	     soc_uart_user_ifc_uart_pwXmitEnableBitCount_whas ;

  // register soc_uart_user_ifc_uart_rXmitCellCount
  assign soc_uart_user_ifc_uart_rXmitCellCount_D_IN =
	     soc_uart_user_ifc_uart_pwXmitCellCountReset_whas ?
	       4'd0 :
	       x__h37182 ;
  assign soc_uart_user_ifc_uart_rXmitCellCount_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // register soc_uart_user_ifc_uart_rXmitDataOut
  always@(MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_1 or
	  soc_uart_user_ifc_uart_vrXmitBuffer_0 or
	  MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_2 or
	  MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_3)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_1:
	  soc_uart_user_ifc_uart_rXmitDataOut_D_IN =
	      soc_uart_user_ifc_uart_vrXmitBuffer_0;
      MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_2:
	  soc_uart_user_ifc_uart_rXmitDataOut_D_IN = 1'b0;
      MUX_soc_uart_user_ifc_uart_rXmitDataOut_write_1__SEL_3:
	  soc_uart_user_ifc_uart_rXmitDataOut_D_IN = 1'b1;
      default: soc_uart_user_ifc_uart_rXmitDataOut_D_IN =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  assign soc_uart_user_ifc_uart_rXmitDataOut_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ;

  // register soc_uart_user_ifc_uart_rXmitParity
  assign soc_uart_user_ifc_uart_rXmitParity_D_IN =
	     z__h38631 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[7] ;
  assign soc_uart_user_ifc_uart_rXmitParity_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ;

  // register soc_uart_user_ifc_uart_rXmitState
  always@(WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_1 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_2 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_3 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_4 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_5 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_6 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 or
	  MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_7 or
	  WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_1;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_2;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_3;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_4;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_5;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_6;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2:
	  soc_uart_user_ifc_uart_rXmitState_D_IN =
	      MUX_soc_uart_user_ifc_uart_rXmitState_write_1__VAL_7;
      WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit:
	  soc_uart_user_ifc_uart_rXmitState_D_IN = 3'd2;
      default: soc_uart_user_ifc_uart_rXmitState_D_IN =
		   3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_uart_user_ifc_uart_rXmitState_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_for_start_command ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit1_5 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_shift_next_bit ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_0
  assign soc_uart_user_ifc_uart_vrRecvBuffer_0_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_1 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_0_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_1
  assign soc_uart_user_ifc_uart_vrRecvBuffer_1_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_2 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_1_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_2
  assign soc_uart_user_ifc_uart_vrRecvBuffer_2_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_3 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_2_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_3
  assign soc_uart_user_ifc_uart_vrRecvBuffer_3_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_4 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_3_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_4
  assign soc_uart_user_ifc_uart_vrRecvBuffer_4_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_5 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_4_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_5
  assign soc_uart_user_ifc_uart_vrRecvBuffer_5_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_6 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_5_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_6
  assign soc_uart_user_ifc_uart_vrRecvBuffer_6_D_IN =
	     soc_uart_user_ifc_uart_vrRecvBuffer_7 ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_6_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrRecvBuffer_7
  assign soc_uart_user_ifc_uart_vrRecvBuffer_7_D_IN =
	     soc_uart_user_ifc_uart_rRecvData ;
  assign soc_uart_user_ifc_uart_vrRecvBuffer_7_EN =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_0
  assign soc_uart_user_ifc_uart_vrXmitBuffer_0_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[0] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_1 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_0_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_1
  assign soc_uart_user_ifc_uart_vrXmitBuffer_1_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[1] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_2 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_1_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_2
  assign soc_uart_user_ifc_uart_vrXmitBuffer_2_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[2] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_3 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_2_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_3
  assign soc_uart_user_ifc_uart_vrXmitBuffer_3_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[3] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_4 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_3_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_4
  assign soc_uart_user_ifc_uart_vrXmitBuffer_4_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[4] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_5 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_4_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_5
  assign soc_uart_user_ifc_uart_vrXmitBuffer_5_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[5] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_6 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_5_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_6
  assign soc_uart_user_ifc_uart_vrXmitBuffer_6_D_IN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ?
	       soc_uart_user_ifc_uart_fifoXmit_D_OUT[6] :
	       soc_uart_user_ifc_uart_vrXmitBuffer_7 ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_6_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // register soc_uart_user_ifc_uart_vrXmitBuffer_7
  assign soc_uart_user_ifc_uart_vrXmitBuffer_7_D_IN =
	     !WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     soc_uart_user_ifc_uart_fifoXmit_D_OUT[7] ;
  assign soc_uart_user_ifc_uart_vrXmitBuffer_7_EN =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_shift ;

  // submodule soc_clint_s_xactor_f_rd_addr
  assign soc_clint_s_xactor_f_rd_addr_D_IN =
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_D_OUT ;
  assign soc_clint_s_xactor_f_rd_addr_ENQ =
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_rd_addr_FULL_N ;
  assign soc_clint_s_xactor_f_rd_addr_DEQ =
	     CAN_FIRE_RL_soc_clint_axi_read_transaction ;
  assign soc_clint_s_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_clint_s_xactor_f_rd_data
  assign soc_clint_s_xactor_f_rd_data_D_IN =
	     { (soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] == 16'h0 ||
		soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] >= 16'h4000 &&
		soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] <= 16'd16391 ||
		soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] >= 16'hBFF8 &&
		soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] <= 16'd49151) ?
		 2'd0 :
		 2'd2,
	       IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078 } ;
  assign soc_clint_s_xactor_f_rd_data_ENQ =
	     CAN_FIRE_RL_soc_clint_axi_read_transaction ;
  assign soc_clint_s_xactor_f_rd_data_DEQ =
	     soc_fabric_xactors_to_slaves_3_f_rd_data_FULL_N &&
	     soc_clint_s_xactor_f_rd_data_EMPTY_N ;
  assign soc_clint_s_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule soc_clint_s_xactor_f_wr_addr
  assign soc_clint_s_xactor_f_wr_addr_D_IN =
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_D_OUT ;
  assign soc_clint_s_xactor_f_wr_addr_ENQ =
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_addr_FULL_N ;
  assign soc_clint_s_xactor_f_wr_addr_DEQ =
	     CAN_FIRE_RL_soc_clint_axi_write_transaction ;
  assign soc_clint_s_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_clint_s_xactor_f_wr_data
  assign soc_clint_s_xactor_f_wr_data_D_IN =
	     soc_fabric_xactors_to_slaves_3_f_wr_data_D_OUT ;
  assign soc_clint_s_xactor_f_wr_data_ENQ =
	     soc_fabric_xactors_to_slaves_3_f_wr_data_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_data_FULL_N ;
  assign soc_clint_s_xactor_f_wr_data_DEQ =
	     CAN_FIRE_RL_soc_clint_axi_write_transaction ;
  assign soc_clint_s_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule soc_clint_s_xactor_f_wr_resp
  assign soc_clint_s_xactor_f_wr_resp_D_IN =
	     (soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] == 16'h0 ||
	      soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] >= 16'h4000 &&
	      soc_clint_s_xactor_f_wr_addr_D_OUT[20:5] <= 16'd16391) ?
	       2'd0 :
	       2'd2 ;
  assign soc_clint_s_xactor_f_wr_resp_ENQ =
	     CAN_FIRE_RL_soc_clint_axi_write_transaction ;
  assign soc_clint_s_xactor_f_wr_resp_DEQ =
	     soc_fabric_xactors_to_slaves_3_f_wr_resp_FULL_N &&
	     soc_clint_s_xactor_f_wr_resp_EMPTY_N ;
  assign soc_clint_s_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_eclass
  assign soc_eclass_master_d_m_arready_arready =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_FULL_N ;
  assign soc_eclass_master_d_m_awready_awready =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_FULL_N ;
  assign soc_eclass_master_d_m_bvalid_bresp =
	     soc_fabric_xactors_from_masters_1_f_wr_resp_D_OUT ;
  assign soc_eclass_master_d_m_bvalid_bvalid =
	     soc_fabric_xactors_from_masters_1_f_wr_resp_EMPTY_N ;
  assign soc_eclass_master_d_m_rvalid_rdata =
	     soc_fabric_xactors_from_masters_1_f_rd_data_D_OUT[63:0] ;
  assign soc_eclass_master_d_m_rvalid_rresp =
	     soc_fabric_xactors_from_masters_1_f_rd_data_D_OUT[65:64] ;
  assign soc_eclass_master_d_m_rvalid_rvalid =
	     soc_fabric_xactors_from_masters_1_f_rd_data_EMPTY_N ;
  assign soc_eclass_master_d_m_wready_wready =
	     soc_fabric_xactors_from_masters_1_f_wr_data_FULL_N ;
  assign soc_eclass_master_i_m_arready_arready =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_FULL_N ;
  assign soc_eclass_master_i_m_awready_awready =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_FULL_N ;
  assign soc_eclass_master_i_m_bvalid_bresp =
	     soc_fabric_xactors_from_masters_2_f_wr_resp_D_OUT ;
  assign soc_eclass_master_i_m_bvalid_bvalid =
	     soc_fabric_xactors_from_masters_2_f_wr_resp_EMPTY_N ;
  assign soc_eclass_master_i_m_rvalid_rdata =
	     soc_fabric_xactors_from_masters_2_f_rd_data_D_OUT[63:0] ;
  assign soc_eclass_master_i_m_rvalid_rresp =
	     soc_fabric_xactors_from_masters_2_f_rd_data_D_OUT[65:64] ;
  assign soc_eclass_master_i_m_rvalid_rvalid =
	     soc_fabric_xactors_from_masters_2_f_rd_data_EMPTY_N ;
  assign soc_eclass_master_i_m_wready_wready =
	     soc_fabric_xactors_from_masters_2_f_wr_data_FULL_N ;
  assign soc_eclass_sb_clint_msip_put = soc_clint_clint_msip ;
  assign soc_eclass_sb_clint_mtime_put = soc_clint_clint_rgmtime ;
  assign soc_eclass_sb_clint_mtip_put = soc_clint_clint_mtip ;
  assign soc_eclass_sb_ext_interrupt_put = 1'b0 ;
  assign soc_eclass_EN_sb_clint_msip_put = 1'd1 ;
  assign soc_eclass_EN_sb_clint_mtip_put = 1'd1 ;
  assign soc_eclass_EN_sb_clint_mtime_put = 1'd1 ;
  assign soc_eclass_EN_sb_ext_interrupt_put = 1'b0 ;
  assign soc_eclass_EN_io_dump_get = 1'b0 ;

  // submodule soc_err_slave_s_xactor_f_rd_addr
  assign soc_err_slave_s_xactor_f_rd_addr_D_IN =
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_D_OUT ;
  assign soc_err_slave_s_xactor_f_rd_addr_ENQ =
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_rd_addr_FULL_N ;
  assign soc_err_slave_s_xactor_f_rd_addr_DEQ =
	     CAN_FIRE_RL_soc_err_slave_receive_read_request ;
  assign soc_err_slave_s_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_err_slave_s_xactor_f_rd_data
  assign soc_err_slave_s_xactor_f_rd_data_D_IN = 66'h30000000000000000 ;
  assign soc_err_slave_s_xactor_f_rd_data_ENQ =
	     CAN_FIRE_RL_soc_err_slave_receive_read_request ;
  assign soc_err_slave_s_xactor_f_rd_data_DEQ =
	     soc_fabric_xactors_to_slaves_5_f_rd_data_FULL_N &&
	     soc_err_slave_s_xactor_f_rd_data_EMPTY_N ;
  assign soc_err_slave_s_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule soc_err_slave_s_xactor_f_wr_addr
  assign soc_err_slave_s_xactor_f_wr_addr_D_IN =
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_D_OUT ;
  assign soc_err_slave_s_xactor_f_wr_addr_ENQ =
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_addr_FULL_N ;
  assign soc_err_slave_s_xactor_f_wr_addr_DEQ =
	     CAN_FIRE_RL_soc_err_slave_receive_write_request ;
  assign soc_err_slave_s_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_err_slave_s_xactor_f_wr_data
  assign soc_err_slave_s_xactor_f_wr_data_D_IN =
	     soc_fabric_xactors_to_slaves_5_f_wr_data_D_OUT ;
  assign soc_err_slave_s_xactor_f_wr_data_ENQ =
	     soc_fabric_xactors_to_slaves_5_f_wr_data_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_data_FULL_N ;
  assign soc_err_slave_s_xactor_f_wr_data_DEQ =
	     CAN_FIRE_RL_soc_err_slave_receive_write_request ;
  assign soc_err_slave_s_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule soc_err_slave_s_xactor_f_wr_resp
  assign soc_err_slave_s_xactor_f_wr_resp_D_IN = 2'd3 ;
  assign soc_err_slave_s_xactor_f_wr_resp_ENQ =
	     CAN_FIRE_RL_soc_err_slave_receive_write_request ;
  assign soc_err_slave_s_xactor_f_wr_resp_DEQ =
	     soc_fabric_xactors_to_slaves_5_f_wr_resp_FULL_N &&
	     soc_err_slave_s_xactor_f_wr_resp_EMPTY_N ;
  assign soc_err_slave_s_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_err_user_0
  assign soc_fabric_v_f_rd_err_user_0_ENQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_0_DEQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_err_user_1
  assign soc_fabric_v_f_rd_err_user_1_ENQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_1_DEQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_err_user_2
  assign soc_fabric_v_f_rd_err_user_2_ENQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_2_DEQ = 1'b0 ;
  assign soc_fabric_v_f_rd_err_user_2_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_0
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave:
	  soc_fabric_v_f_rd_mis_0_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6:
	  soc_fabric_v_f_rd_mis_0_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12:
	  soc_fabric_v_f_rd_mis_0_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_0_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_0_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 ;
  assign soc_fabric_v_f_rd_mis_0_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master ;
  assign soc_fabric_v_f_rd_mis_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_1
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1:
	  soc_fabric_v_f_rd_mis_1_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7:
	  soc_fabric_v_f_rd_mis_1_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13:
	  soc_fabric_v_f_rd_mis_1_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_1_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_1_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 ;
  assign soc_fabric_v_f_rd_mis_1_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 ;
  assign soc_fabric_v_f_rd_mis_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_2
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2:
	  soc_fabric_v_f_rd_mis_2_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8:
	  soc_fabric_v_f_rd_mis_2_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14:
	  soc_fabric_v_f_rd_mis_2_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_2_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_2_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 ;
  assign soc_fabric_v_f_rd_mis_2_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 ;
  assign soc_fabric_v_f_rd_mis_2_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_3
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3:
	  soc_fabric_v_f_rd_mis_3_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9:
	  soc_fabric_v_f_rd_mis_3_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15:
	  soc_fabric_v_f_rd_mis_3_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_3_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_3_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 ;
  assign soc_fabric_v_f_rd_mis_3_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 ;
  assign soc_fabric_v_f_rd_mis_3_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_4
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4:
	  soc_fabric_v_f_rd_mis_4_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10:
	  soc_fabric_v_f_rd_mis_4_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16:
	  soc_fabric_v_f_rd_mis_4_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_4_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_4_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 ;
  assign soc_fabric_v_f_rd_mis_4_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 ;
  assign soc_fabric_v_f_rd_mis_4_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_mis_5
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5:
	  soc_fabric_v_f_rd_mis_5_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11:
	  soc_fabric_v_f_rd_mis_5_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17:
	  soc_fabric_v_f_rd_mis_5_D_IN = 2'd2;
      default: soc_fabric_v_f_rd_mis_5_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_mis_5_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 ;
  assign soc_fabric_v_f_rd_mis_5_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 ;
  assign soc_fabric_v_f_rd_mis_5_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_sjs_0
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5:
	  soc_fabric_v_f_rd_sjs_0_D_IN = 3'd5;
      default: soc_fabric_v_f_rd_sjs_0_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_sjs_0_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ;
  assign soc_fabric_v_f_rd_sjs_0_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master ;
  assign soc_fabric_v_f_rd_sjs_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_sjs_1
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11:
	  soc_fabric_v_f_rd_sjs_1_D_IN = 3'd5;
      default: soc_fabric_v_f_rd_sjs_1_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_sjs_1_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 ;
  assign soc_fabric_v_f_rd_sjs_1_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 ;
  assign soc_fabric_v_f_rd_sjs_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_rd_sjs_2
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17:
	  soc_fabric_v_f_rd_sjs_2_D_IN = 3'd5;
      default: soc_fabric_v_f_rd_sjs_2_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_rd_sjs_2_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 ;
  assign soc_fabric_v_f_rd_sjs_2_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 ;
  assign soc_fabric_v_f_rd_sjs_2_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_err_user_0
  assign soc_fabric_v_f_wr_err_user_0_ENQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_0_DEQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_err_user_1
  assign soc_fabric_v_f_wr_err_user_1_ENQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_1_DEQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_err_user_2
  assign soc_fabric_v_f_wr_err_user_2_ENQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_2_DEQ = 1'b0 ;
  assign soc_fabric_v_f_wr_err_user_2_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_0
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave:
	  soc_fabric_v_f_wr_mis_0_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6:
	  soc_fabric_v_f_wr_mis_0_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12:
	  soc_fabric_v_f_wr_mis_0_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_0_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_0_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ;
  assign soc_fabric_v_f_wr_mis_0_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master ;
  assign soc_fabric_v_f_wr_mis_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_1
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1:
	  soc_fabric_v_f_wr_mis_1_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7:
	  soc_fabric_v_f_wr_mis_1_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13:
	  soc_fabric_v_f_wr_mis_1_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_1_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_1_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ;
  assign soc_fabric_v_f_wr_mis_1_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 ;
  assign soc_fabric_v_f_wr_mis_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_2
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2:
	  soc_fabric_v_f_wr_mis_2_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8:
	  soc_fabric_v_f_wr_mis_2_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14:
	  soc_fabric_v_f_wr_mis_2_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_2_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_2_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ;
  assign soc_fabric_v_f_wr_mis_2_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 ;
  assign soc_fabric_v_f_wr_mis_2_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_3
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3:
	  soc_fabric_v_f_wr_mis_3_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9:
	  soc_fabric_v_f_wr_mis_3_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15:
	  soc_fabric_v_f_wr_mis_3_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_3_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_3_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ;
  assign soc_fabric_v_f_wr_mis_3_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 ;
  assign soc_fabric_v_f_wr_mis_3_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_4
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4:
	  soc_fabric_v_f_wr_mis_4_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10:
	  soc_fabric_v_f_wr_mis_4_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16:
	  soc_fabric_v_f_wr_mis_4_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_4_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_4_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ;
  assign soc_fabric_v_f_wr_mis_4_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 ;
  assign soc_fabric_v_f_wr_mis_4_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_mis_5
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5:
	  soc_fabric_v_f_wr_mis_5_D_IN = 2'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11:
	  soc_fabric_v_f_wr_mis_5_D_IN = 2'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17:
	  soc_fabric_v_f_wr_mis_5_D_IN = 2'd2;
      default: soc_fabric_v_f_wr_mis_5_D_IN = 2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_mis_5_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ;
  assign soc_fabric_v_f_wr_mis_5_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 ;
  assign soc_fabric_v_f_wr_mis_5_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_sjs_0
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5:
	  soc_fabric_v_f_wr_sjs_0_D_IN = 3'd5;
      default: soc_fabric_v_f_wr_sjs_0_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_sjs_0_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ;
  assign soc_fabric_v_f_wr_sjs_0_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master ;
  assign soc_fabric_v_f_wr_sjs_0_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_sjs_1
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11:
	  soc_fabric_v_f_wr_sjs_1_D_IN = 3'd5;
      default: soc_fabric_v_f_wr_sjs_1_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_sjs_1_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ;
  assign soc_fabric_v_f_wr_sjs_1_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 ;
  assign soc_fabric_v_f_wr_sjs_1_CLR = 1'b0 ;

  // submodule soc_fabric_v_f_wr_sjs_2
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd0;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd1;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd2;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd3;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd4;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17:
	  soc_fabric_v_f_wr_sjs_2_D_IN = 3'd5;
      default: soc_fabric_v_f_wr_sjs_2_D_IN = 3'b010 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_v_f_wr_sjs_2_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ;
  assign soc_fabric_v_f_wr_sjs_2_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 ;
  assign soc_fabric_v_f_wr_sjs_2_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_0_f_rd_addr
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_D_IN =
	     { soc_signature_master_araddr,
	       soc_signature_master_arprot,
	       soc_signature_master_arsize } ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_ENQ =
	     soc_signature_master_arvalid &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_0_f_rd_data
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master or
	  soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 or
	  soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 or
	  soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 or
	  soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 or
	  soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 or
	  soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5:
	  soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT;
      default: soc_fabric_xactors_from_masters_0_f_rd_data_D_IN =
		   66'h2AAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_0_f_rd_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_data_DEQ =
	     soc_signature_master_rready &&
	     soc_fabric_xactors_from_masters_0_f_rd_data_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_0_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_0_f_wr_addr
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_D_IN =
	     { soc_signature_master_awaddr,
	       soc_signature_master_awprot,
	       soc_signature_master_awsize } ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_ENQ =
	     soc_signature_master_awvalid &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_0_f_wr_data
  assign soc_fabric_xactors_from_masters_0_f_wr_data_D_IN =
	     { soc_signature_master_wdata, soc_signature_master_wstrb } ;
  assign soc_fabric_xactors_from_masters_0_f_wr_data_ENQ =
	     soc_signature_master_wvalid &&
	     soc_fabric_xactors_from_masters_0_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_from_masters_0_f_wr_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ;
  assign soc_fabric_xactors_from_masters_0_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_0_f_wr_resp
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master or
	  soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 or
	  soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 or
	  soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 or
	  soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 or
	  soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 or
	  soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5:
	  soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT;
      default: soc_fabric_xactors_from_masters_0_f_wr_resp_D_IN =
		   2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_0_f_wr_resp_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_resp_DEQ =
	     soc_signature_master_bready &&
	     soc_fabric_xactors_from_masters_0_f_wr_resp_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_0_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_1_f_rd_addr
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_D_IN =
	     { soc_eclass_master_d_araddr,
	       soc_eclass_master_d_arprot,
	       soc_eclass_master_d_arsize } ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_ENQ =
	     soc_eclass_master_d_arvalid &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_1_f_rd_data
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 or
	  soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 or
	  soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 or
	  soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 or
	  soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 or
	  soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 or
	  soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11:
	  soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT;
      default: soc_fabric_xactors_from_masters_1_f_rd_data_D_IN =
		   66'h2AAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_1_f_rd_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_data_DEQ =
	     soc_eclass_master_d_rready &&
	     soc_fabric_xactors_from_masters_1_f_rd_data_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_1_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_1_f_wr_addr
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_D_IN =
	     { soc_eclass_master_d_awaddr,
	       soc_eclass_master_d_awprot,
	       soc_eclass_master_d_awsize } ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_ENQ =
	     soc_eclass_master_d_awvalid &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_1_f_wr_data
  assign soc_fabric_xactors_from_masters_1_f_wr_data_D_IN =
	     { soc_eclass_master_d_wdata, soc_eclass_master_d_wstrb } ;
  assign soc_fabric_xactors_from_masters_1_f_wr_data_ENQ =
	     soc_eclass_master_d_wvalid &&
	     soc_fabric_xactors_from_masters_1_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_from_masters_1_f_wr_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_1_f_wr_resp
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 or
	  soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 or
	  soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 or
	  soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 or
	  soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 or
	  soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 or
	  soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11:
	  soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT;
      default: soc_fabric_xactors_from_masters_1_f_wr_resp_D_IN =
		   2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_1_f_wr_resp_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_resp_DEQ =
	     soc_eclass_master_d_bready &&
	     soc_fabric_xactors_from_masters_1_f_wr_resp_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_1_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_2_f_rd_addr
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_D_IN =
	     { soc_eclass_master_i_araddr,
	       soc_eclass_master_i_arprot,
	       soc_eclass_master_i_arsize } ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_ENQ =
	     soc_eclass_master_i_arvalid &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_2_f_rd_data
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 or
	  soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 or
	  soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 or
	  soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 or
	  soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 or
	  soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 or
	  soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_rd_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17:
	  soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_rd_data_D_OUT;
      default: soc_fabric_xactors_from_masters_2_f_rd_data_D_IN =
		   66'h2AAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_2_f_rd_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_data_DEQ =
	     soc_eclass_master_i_rready &&
	     soc_fabric_xactors_from_masters_2_f_rd_data_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_2_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_2_f_wr_addr
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_D_IN =
	     { soc_eclass_master_i_awaddr,
	       soc_eclass_master_i_awprot,
	       soc_eclass_master_i_awsize } ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_ENQ =
	     soc_eclass_master_i_awvalid &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_2_f_wr_data
  assign soc_fabric_xactors_from_masters_2_f_wr_data_D_IN =
	     { soc_eclass_master_i_wdata, soc_eclass_master_i_wstrb } ;
  assign soc_fabric_xactors_from_masters_2_f_wr_data_ENQ =
	     soc_eclass_master_i_wvalid &&
	     soc_fabric_xactors_from_masters_2_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_from_masters_2_f_wr_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_from_masters_2_f_wr_resp
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 or
	  soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 or
	  soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 or
	  soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 or
	  soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 or
	  soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 or
	  soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_0_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_1_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_2_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_3_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_4_f_wr_resp_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17:
	  soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
	      soc_fabric_xactors_to_slaves_5_f_wr_resp_D_OUT;
      default: soc_fabric_xactors_from_masters_2_f_wr_resp_D_IN =
		   2'b10 /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_from_masters_2_f_wr_resp_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_resp_DEQ =
	     soc_eclass_master_i_bready &&
	     soc_fabric_xactors_from_masters_2_f_wr_resp_EMPTY_N ;
  assign soc_fabric_xactors_from_masters_2_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_0_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave:
	  soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6:
	  soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12:
	  soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_0_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_0_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_to_slaves_0_f_rd_addr_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_0_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_0_f_rd_data
  assign soc_fabric_xactors_to_slaves_0_f_rd_data_D_IN = 66'h0 ;
  assign soc_fabric_xactors_to_slaves_0_f_rd_data_ENQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_0_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master ;
  assign soc_fabric_xactors_to_slaves_0_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave:
	  soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6:
	  soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12:
	  soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_0_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_0_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_addr_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave:
	  soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6:
	  soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12:
	  soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_0_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_0_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_12 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_data_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_0_f_wr_resp
  assign soc_fabric_xactors_to_slaves_0_f_wr_resp_D_IN = 2'h0 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_resp_ENQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_12 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_6 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master ;
  assign soc_fabric_xactors_to_slaves_0_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_1_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1:
	  soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7:
	  soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13:
	  soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_1_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_1_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_13 ;
  assign soc_fabric_xactors_to_slaves_1_f_rd_addr_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_1_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_1_f_rd_data
  assign soc_fabric_xactors_to_slaves_1_f_rd_data_D_IN = 66'h0 ;
  assign soc_fabric_xactors_to_slaves_1_f_rd_data_ENQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_1_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_1 ;
  assign soc_fabric_xactors_to_slaves_1_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1:
	  soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7:
	  soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13:
	  soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_1_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_1_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_addr_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1:
	  soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7:
	  soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13:
	  soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_1_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_1_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_1 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_13 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_data_DEQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_1_f_wr_resp
  assign soc_fabric_xactors_to_slaves_1_f_wr_resp_D_IN = 2'h0 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_resp_ENQ = 1'b0 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_13 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_7 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_1 ;
  assign soc_fabric_xactors_to_slaves_1_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_2_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2:
	  soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8:
	  soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14:
	  soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_2_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_2_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_14 ;
  assign soc_fabric_xactors_to_slaves_2_f_rd_addr_DEQ =
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_2_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_2_f_rd_data
  assign soc_fabric_xactors_to_slaves_2_f_rd_data_D_IN =
	     soc_uart_s_xactor_f_rd_data_D_OUT ;
  assign soc_fabric_xactors_to_slaves_2_f_rd_data_ENQ =
	     soc_uart_s_xactor_f_rd_data_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_rd_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_2_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_2 ;
  assign soc_fabric_xactors_to_slaves_2_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2:
	  soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8:
	  soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14:
	  soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_2_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_2_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_addr_DEQ =
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2:
	  soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8:
	  soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14:
	  soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_2_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_2_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_2 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_14 ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_data_DEQ =
	     soc_fabric_xactors_to_slaves_2_f_wr_data_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_2_f_wr_resp
  assign soc_fabric_xactors_to_slaves_2_f_wr_resp_D_IN =
	     soc_uart_s_xactor_f_wr_resp_D_OUT ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_resp_ENQ =
	     soc_uart_s_xactor_f_wr_resp_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_2_f_wr_resp_FULL_N ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_14 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_8 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_2 ;
  assign soc_fabric_xactors_to_slaves_2_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_3_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3:
	  soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9:
	  soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15:
	  soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_3_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_3_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_15 ;
  assign soc_fabric_xactors_to_slaves_3_f_rd_addr_DEQ =
	     soc_fabric_xactors_to_slaves_3_f_rd_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_3_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_3_f_rd_data
  assign soc_fabric_xactors_to_slaves_3_f_rd_data_D_IN =
	     soc_clint_s_xactor_f_rd_data_D_OUT ;
  assign soc_fabric_xactors_to_slaves_3_f_rd_data_ENQ =
	     soc_clint_s_xactor_f_rd_data_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_rd_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_3_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_3 ;
  assign soc_fabric_xactors_to_slaves_3_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3:
	  soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9:
	  soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15:
	  soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_3_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_3_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_addr_DEQ =
	     soc_fabric_xactors_to_slaves_3_f_wr_addr_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3:
	  soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9:
	  soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15:
	  soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_3_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_3_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_3 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_15 ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_data_DEQ =
	     soc_fabric_xactors_to_slaves_3_f_wr_data_EMPTY_N &&
	     soc_clint_s_xactor_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_3_f_wr_resp
  assign soc_fabric_xactors_to_slaves_3_f_wr_resp_D_IN =
	     soc_clint_s_xactor_f_wr_resp_D_OUT ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_resp_ENQ =
	     soc_clint_s_xactor_f_wr_resp_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_3_f_wr_resp_FULL_N ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_15 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_9 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_3 ;
  assign soc_fabric_xactors_to_slaves_3_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_4_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4:
	  soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10:
	  soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16:
	  soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_4_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_4_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_16 ;
  assign soc_fabric_xactors_to_slaves_4_f_rd_addr_DEQ =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_EMPTY_N &&
	     soc_signature_slave_arready ;
  assign soc_fabric_xactors_to_slaves_4_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_4_f_rd_data
  assign soc_fabric_xactors_to_slaves_4_f_rd_data_D_IN =
	     { soc_signature_slave_rresp, soc_signature_slave_rdata } ;
  assign soc_fabric_xactors_to_slaves_4_f_rd_data_ENQ =
	     soc_signature_slave_rvalid &&
	     soc_fabric_xactors_to_slaves_4_f_rd_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_4_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_4 ;
  assign soc_fabric_xactors_to_slaves_4_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4:
	  soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10:
	  soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16:
	  soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_4_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_4_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_addr_DEQ =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_EMPTY_N &&
	     soc_signature_slave_awready ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4:
	  soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10:
	  soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16:
	  soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_4_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_4_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_4 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_16 ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_data_DEQ =
	     soc_fabric_xactors_to_slaves_4_f_wr_data_EMPTY_N &&
	     soc_signature_slave_wready ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_4_f_wr_resp
  assign soc_fabric_xactors_to_slaves_4_f_wr_resp_D_IN =
	     soc_signature_slave_bresp ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_resp_ENQ =
	     soc_signature_slave_bvalid &&
	     soc_fabric_xactors_to_slaves_4_f_wr_resp_FULL_N ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_16 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_10 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_4 ;
  assign soc_fabric_xactors_to_slaves_4_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_5_f_rd_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 or
	  soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 or
	  soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 or
	  soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5:
	  soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11:
	  soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17:
	  soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_5_f_rd_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_5_f_rd_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_xaction_master_to_slave_17 ;
  assign soc_fabric_xactors_to_slaves_5_f_rd_addr_DEQ =
	     soc_fabric_xactors_to_slaves_5_f_rd_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_rd_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_5_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_5_f_rd_data
  assign soc_fabric_xactors_to_slaves_5_f_rd_data_D_IN =
	     soc_err_slave_s_xactor_f_rd_data_D_OUT ;
  assign soc_fabric_xactors_to_slaves_5_f_rd_data_ENQ =
	     soc_err_slave_s_xactor_f_rd_data_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_rd_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_5_f_rd_data_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_rd_resp_slave_to_master_5 ;
  assign soc_fabric_xactors_to_slaves_5_f_rd_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_addr
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 or
	  soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 or
	  soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 or
	  soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5:
	  soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11:
	  soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17:
	  soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT;
      default: soc_fabric_xactors_to_slaves_5_f_wr_addr_D_IN =
		   37'h0AAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_5_f_wr_addr_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_addr_DEQ =
	     soc_fabric_xactors_to_slaves_5_f_wr_addr_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_addr_FULL_N ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_data
  always@(WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 or
	  soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 or
	  soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT or
	  WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 or
	  soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5:
	  soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_0_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11:
	  soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_1_f_wr_data_D_OUT;
      WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17:
	  soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN =
	      soc_fabric_xactors_from_masters_2_f_wr_data_D_OUT;
      default: soc_fabric_xactors_to_slaves_5_f_wr_data_D_IN =
		   72'hAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign soc_fabric_xactors_to_slaves_5_f_wr_data_ENQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_5 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_xaction_master_to_slave_17 ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_data_DEQ =
	     soc_fabric_xactors_to_slaves_5_f_wr_data_EMPTY_N &&
	     soc_err_slave_s_xactor_f_wr_data_FULL_N ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_data_CLR = 1'b0 ;

  // submodule soc_fabric_xactors_to_slaves_5_f_wr_resp
  assign soc_fabric_xactors_to_slaves_5_f_wr_resp_D_IN =
	     soc_err_slave_s_xactor_f_wr_resp_D_OUT ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_resp_ENQ =
	     soc_err_slave_s_xactor_f_wr_resp_EMPTY_N &&
	     soc_fabric_xactors_to_slaves_5_f_wr_resp_FULL_N ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_resp_DEQ =
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_17 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_11 ||
	     WILL_FIRE_RL_soc_fabric_rl_wr_resp_slave_to_master_5 ;
  assign soc_fabric_xactors_to_slaves_5_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_signature
  assign soc_signature_master_m_arready_arready =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_FULL_N ;
  assign soc_signature_master_m_awready_awready =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_FULL_N ;
  assign soc_signature_master_m_bvalid_bresp =
	     soc_fabric_xactors_from_masters_0_f_wr_resp_D_OUT ;
  assign soc_signature_master_m_bvalid_bvalid =
	     soc_fabric_xactors_from_masters_0_f_wr_resp_EMPTY_N ;
  assign soc_signature_master_m_rvalid_rdata =
	     soc_fabric_xactors_from_masters_0_f_rd_data_D_OUT[63:0] ;
  assign soc_signature_master_m_rvalid_rresp =
	     soc_fabric_xactors_from_masters_0_f_rd_data_D_OUT[65:64] ;
  assign soc_signature_master_m_rvalid_rvalid =
	     soc_fabric_xactors_from_masters_0_f_rd_data_EMPTY_N ;
  assign soc_signature_master_m_wready_wready =
	     soc_fabric_xactors_from_masters_0_f_wr_data_FULL_N ;
  assign soc_signature_slave_m_arvalid_araddr =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_D_OUT[36:5] ;
  assign soc_signature_slave_m_arvalid_arprot =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_D_OUT[4:2] ;
  assign soc_signature_slave_m_arvalid_arsize =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_D_OUT[1:0] ;
  assign soc_signature_slave_m_arvalid_arvalid =
	     soc_fabric_xactors_to_slaves_4_f_rd_addr_EMPTY_N ;
  assign soc_signature_slave_m_awvalid_awaddr =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_D_OUT[36:5] ;
  assign soc_signature_slave_m_awvalid_awprot =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_D_OUT[4:2] ;
  assign soc_signature_slave_m_awvalid_awsize =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_D_OUT[1:0] ;
  assign soc_signature_slave_m_awvalid_awvalid =
	     soc_fabric_xactors_to_slaves_4_f_wr_addr_EMPTY_N ;
  assign soc_signature_slave_m_bready_bready =
	     soc_fabric_xactors_to_slaves_4_f_wr_resp_FULL_N ;
  assign soc_signature_slave_m_rready_rready =
	     soc_fabric_xactors_to_slaves_4_f_rd_data_FULL_N ;
  assign soc_signature_slave_m_wvalid_wdata =
	     soc_fabric_xactors_to_slaves_4_f_wr_data_D_OUT[71:8] ;
  assign soc_signature_slave_m_wvalid_wstrb =
	     soc_fabric_xactors_to_slaves_4_f_wr_data_D_OUT[7:0] ;
  assign soc_signature_slave_m_wvalid_wvalid =
	     soc_fabric_xactors_to_slaves_4_f_wr_data_EMPTY_N ;

  // submodule soc_uart_s_xactor_f_rd_addr
  assign soc_uart_s_xactor_f_rd_addr_D_IN =
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_D_OUT ;
  assign soc_uart_s_xactor_f_rd_addr_ENQ =
	     soc_fabric_xactors_to_slaves_2_f_rd_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_rd_addr_FULL_N ;
  assign soc_uart_s_xactor_f_rd_addr_DEQ =
	     CAN_FIRE_RL_soc_uart_capture_read_request ;
  assign soc_uart_s_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule soc_uart_s_xactor_f_rd_data
  assign soc_uart_s_xactor_f_rd_data_D_IN =
	     { (soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'hC &&
		soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0 ||
		soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'h8 &&
		soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0 ||
		soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'h0 &&
		soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd1) ?
		 2'd0 :
		 2'd2,
	       IF_soc_uart_s_xactor_f_rd_addr_first__39_BITS__ETC___d971 } ;
  assign soc_uart_s_xactor_f_rd_data_ENQ =
	     CAN_FIRE_RL_soc_uart_capture_read_request ;
  assign soc_uart_s_xactor_f_rd_data_DEQ =
	     soc_fabric_xactors_to_slaves_2_f_rd_data_FULL_N &&
	     soc_uart_s_xactor_f_rd_data_EMPTY_N ;
  assign soc_uart_s_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule soc_uart_s_xactor_f_wr_addr
  assign soc_uart_s_xactor_f_wr_addr_D_IN =
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_D_OUT ;
  assign soc_uart_s_xactor_f_wr_addr_ENQ =
	     soc_fabric_xactors_to_slaves_2_f_wr_addr_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_addr_FULL_N ;
  assign soc_uart_s_xactor_f_wr_addr_DEQ =
	     CAN_FIRE_RL_soc_uart_capture_write_request ;
  assign soc_uart_s_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule soc_uart_s_xactor_f_wr_data
  assign soc_uart_s_xactor_f_wr_data_D_IN =
	     soc_fabric_xactors_to_slaves_2_f_wr_data_D_OUT ;
  assign soc_uart_s_xactor_f_wr_data_ENQ =
	     soc_fabric_xactors_to_slaves_2_f_wr_data_EMPTY_N &&
	     soc_uart_s_xactor_f_wr_data_FULL_N ;
  assign soc_uart_s_xactor_f_wr_data_DEQ =
	     CAN_FIRE_RL_soc_uart_capture_write_request ;
  assign soc_uart_s_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule soc_uart_s_xactor_f_wr_resp
  assign soc_uart_s_xactor_f_wr_resp_D_IN =
	     (soc_uart_s_xactor_f_wr_addr_D_OUT[8:5] == 4'h4 &&
	      soc_uart_s_xactor_f_wr_addr_D_OUT[1:0] == 2'd0 ||
	      soc_uart_s_xactor_f_wr_addr_D_OUT[8:5] == 4'h0 &&
	      soc_uart_s_xactor_f_wr_addr_D_OUT[1:0] == 2'd1) ?
	       2'd0 :
	       2'd2 ;
  assign soc_uart_s_xactor_f_wr_resp_ENQ =
	     CAN_FIRE_RL_soc_uart_capture_write_request ;
  assign soc_uart_s_xactor_f_wr_resp_DEQ =
	     soc_fabric_xactors_to_slaves_2_f_wr_resp_FULL_N &&
	     soc_uart_s_xactor_f_wr_resp_EMPTY_N ;
  assign soc_uart_s_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule soc_uart_user_ifc_uart_baudGen_rBaudCounter
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_A = 16'd1 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_B = 16'h0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_C = 16'h0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_DATA_F = 16'd0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDA =
	     soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_ADDB = 1'b0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETC = 1'b0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_SETF =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;

  // submodule soc_uart_user_ifc_uart_baudGen_rBaudTickCounter
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_A = 3'd1 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_B = 3'h0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_C = 3'h0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_DATA_F = 3'h0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDA =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_baudGen_count_baudtick_16x ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_ADDB = 1'b0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETC = 1'b0 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudTickCounter_SETF = 1'b0 ;

  // submodule soc_uart_user_ifc_uart_fifoRecv
  assign soc_uart_user_ifc_uart_fifoRecv_D_IN =
	     { soc_uart_user_ifc_uart_vrRecvBuffer_7,
	       soc_uart_user_ifc_uart_vrRecvBuffer_6,
	       soc_uart_user_ifc_uart_vrRecvBuffer_5,
	       soc_uart_user_ifc_uart_vrRecvBuffer_4,
	       soc_uart_user_ifc_uart_vrRecvBuffer_3,
	       soc_uart_user_ifc_uart_vrRecvBuffer_2,
	       soc_uart_user_ifc_uart_vrRecvBuffer_1,
	       soc_uart_user_ifc_uart_vrRecvBuffer_0 } ;
  assign soc_uart_user_ifc_uart_fifoRecv_ENQ =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_receive_stop_last_bit ;
  assign soc_uart_user_ifc_uart_fifoRecv_DEQ =
	     soc_uart_user_ifc_uart_fifoRecv_r_deq_whas ;
  assign soc_uart_user_ifc_uart_fifoRecv_CLR = 1'b0 ;

  // submodule soc_uart_user_ifc_uart_fifoXmit
  assign soc_uart_user_ifc_uart_fifoXmit_D_IN =
	     soc_uart_s_xactor_f_wr_data_D_OUT[15:8] ;
  assign soc_uart_user_ifc_uart_fifoXmit_ENQ =
	     soc_uart_user_ifc_uart_fifoXmit_r_enq_whas ;
  assign soc_uart_user_ifc_uart_fifoXmit_DEQ =
	     CAN_FIRE_RL_soc_uart_user_ifc_uart_transmit_buffer_load ;
  assign soc_uart_user_ifc_uart_fifoXmit_CLR = 1'b0 ;

  // remaining internal signals
  assign IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1070 =
	     (soc_clint_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0) ?
	       temp___1__h47250 :
	       temp__h46605 ;
  assign IF_soc_uart_s_xactor_f_rd_addr_first__39_BITS__ETC___d971 =
	     (soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'hC &&
	      soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0) ?
	       a__h41688 :
	       ((soc_uart_s_xactor_f_rd_addr_D_OUT[8:5] == 4'h8 &&
		 soc_uart_s_xactor_f_rd_addr_D_OUT[1:0] == 2'd0) ?
		  a__h41694 :
		  a__h41696) ;
  assign _dor2soc_uart_user_ifc_uart_pwXmitCellCountReset_EN_wset =
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit2 ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_stop_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_parity_bit ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_wait_1_bit_cell_time ||
	     WILL_FIRE_RL_soc_uart_user_ifc_uart_transmit_send_start_bit ;
  assign _theResult___snd__h46661 =
	     (soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] == 16'h0) ?
	       temp___1__h46656 :
	       _theResult___snd__h46728 ;
  assign _theResult___snd__h46728 =
	     (soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] >= 16'h4000 &&
	      soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] <= 16'd16391) ?
	       soc_clint_clint_rgmtimecmp :
	       _theResult___snd__h46795 ;
  assign _theResult___snd__h46795 =
	     (soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] >= 16'hBFF8 &&
	      soc_clint_s_xactor_f_rd_addr_D_OUT[20:5] <= 16'd49151) ?
	       soc_clint_clint_rgmtime :
	       64'd0 ;
  assign a__h41688 = {16{soc_uart_user_ifc_wr_status_wget}} ;
  assign a__h41694 = {8{soc_uart_user_ifc_uart_fifoRecv_D_OUT}} ;
  assign a__h41696 = {4{soc_uart_user_ifc_baud_value}} ;
  assign datamask__h56751 = data__h56748 & mask__h56750 ;
  assign mask__h56750 = mask__h56747 << shift_amt__h56749 ;
  assign notmask__h56752 = ~mask__h56750 ;
  assign shift_amt__h46602 =
	     { soc_clint_s_xactor_f_rd_addr_D_OUT[7:5], 3'd0 } ;
  assign shift_amt__h56749 =
	     { soc_clint_s_xactor_f_wr_addr_D_OUT[7:5], 3'd0 } ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d296 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280) &&
	     !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291 &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d305 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d307 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d310 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293) &&
	     !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d305 &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d307 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d320 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d322 =
	     soc_fabric_xactors_from_masters_0_f_rd_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d325 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d305 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d307) &&
	     !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d320 &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d322 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d327 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280) &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d325 ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d337 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d291 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d293) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d305 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d307) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d320 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d322) ;
  assign soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d339 =
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d266 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d268) &&
	     (soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d278 ||
	      !soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d280) &&
	     soc_fabric_xactors_from_masters_0_f_rd_addr_fi_ETC___d337 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d101 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d63 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d65) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d81 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d83) ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d103 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32) &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d101 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d51 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32) &&
	     !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46 &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d63 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d65 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d68 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48) &&
	     !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d63 &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d65 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d81 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d83 =
	     soc_fabric_xactors_from_masters_0_f_wr_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d86 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d46 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d48) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d63 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d65) &&
	     !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d81 &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d83 ;
  assign soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d88 =
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d14 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d16) &&
	     (soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d30 ||
	      !soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d32) &&
	     soc_fabric_xactors_from_masters_0_f_wr_addr_fi_ETC___d86 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d372 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359) &&
	     !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367 &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d378 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d380 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d383 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369) &&
	     !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d378 &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d380 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d390 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d392 =
	     soc_fabric_xactors_from_masters_1_f_rd_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d395 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d378 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d380) &&
	     !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d390 &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d392 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d397 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359) &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d395 ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d404 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d367 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d369) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d378 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d380) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d390 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d392) ;
  assign soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d406 =
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d348 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d350) &&
	     (soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d357 ||
	      !soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d359) &&
	     soc_fabric_xactors_from_masters_1_f_rd_addr_fi_ETC___d404 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d142 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128) &&
	     !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137 &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d149 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d151 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d154 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139) &&
	     !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d149 &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d151 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d162 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d164 =
	     soc_fabric_xactors_from_masters_1_f_wr_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d167 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d149 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d151) &&
	     !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d162 &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d164 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d169 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128) &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d167 ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d177 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d137 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d139) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d149 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d151) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d162 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d164) ;
  assign soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d179 =
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d115 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d117) &&
	     (soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d126 ||
	      !soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d128) &&
	     soc_fabric_xactors_from_masters_1_f_wr_addr_fi_ETC___d177 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d439 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426) &&
	     !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434 &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d445 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d447 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d450 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436) &&
	     !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d445 &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d447 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d457 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d459 =
	     soc_fabric_xactors_from_masters_2_f_rd_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d462 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d445 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d447) &&
	     !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d457 &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d459 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d464 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426) &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d462 ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d471 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d434 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d436) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d445 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d447) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d457 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d459) ;
  assign soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d473 =
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d415 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d417) &&
	     (soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d424 ||
	      !soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d426) &&
	     soc_fabric_xactors_from_masters_2_f_rd_addr_fi_ETC___d471 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <
	     32'h80000000 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <=
	     32'h8FFFFFFF ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <
	     32'h00001000 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <=
	     32'h00010FFF ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <
	     32'h00011300 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <=
	     32'h00011340 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d218 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204) &&
	     !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213 &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d225 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <
	     32'h02000000 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d227 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <=
	     32'h020BFFFF ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d230 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215) &&
	     !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d225 &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d227 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d238 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <
	     32'h00020000 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d240 =
	     soc_fabric_xactors_from_masters_2_f_wr_addr_D_OUT[36:5] <=
	     32'h0002000C ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d243 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d225 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d227) &&
	     !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d238 &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d240 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d245 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204) &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d243 ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d253 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d213 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d215) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d225 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d227) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d238 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d240) ;
  assign soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d255 =
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d191 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d193) &&
	     (soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d202 ||
	      !soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d204) &&
	     soc_fabric_xactors_from_masters_2_f_wr_addr_fi_ETC___d253 ;
  assign soc_uart_user_ifc_uart_baudGen_rBaudCounter_va_ETC___d802 =
	     soc_uart_user_ifc_uart_baudGen_rBaudCounter_Q_OUT + 16'd1 <
	     soc_uart_user_ifc_baud_value ;
  assign temp___1__h46656 = {64{soc_clint_clint_msip}} ;
  assign temp___1__h47250 = {8{temp__h46605[7:0]}} ;
  assign temp__h46605 = _theResult___snd__h46661 >> shift_amt__h46602 ;
  assign temp__h46821 =
	     {4{IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1070[15:0]}} ;
  assign temp__h56130 =
	     {2{IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1070[31:0]}} ;
  assign x__h33749 = soc_uart_user_ifc_uart_rRecvCellCount + 4'd1 ;
  assign x__h35390 = soc_uart_user_ifc_uart_rRecvBitCount + 4'd1 ;
  assign x__h37182 = soc_uart_user_ifc_uart_rXmitCellCount + 4'd1 ;
  assign x__h37208 = soc_uart_user_ifc_uart_rXmitBitCount + 4'd1 ;
  assign x__h58828 = soc_clint_clint_rgmtimecmp & notmask__h56752 ;
  assign z__h38596 =
	     soc_uart_user_ifc_uart_fifoXmit_D_OUT[0] ^
	     soc_uart_user_ifc_uart_fifoXmit_D_OUT[1] ;
  assign z__h38603 = z__h38596 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[2] ;
  assign z__h38610 = z__h38603 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[3] ;
  assign z__h38617 = z__h38610 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[4] ;
  assign z__h38624 = z__h38617 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[5] ;
  assign z__h38631 = z__h38624 ^ soc_uart_user_ifc_uart_fifoXmit_D_OUT[6] ;
  always@(soc_clint_s_xactor_f_wr_addr_D_OUT or
	  soc_clint_s_xactor_f_wr_data_D_OUT)
  begin
    case (soc_clint_s_xactor_f_wr_addr_D_OUT[1:0])
      2'd0: data__h56748 = {8{soc_clint_s_xactor_f_wr_data_D_OUT[15:8]}};
      2'd1: data__h56748 = {4{soc_clint_s_xactor_f_wr_data_D_OUT[23:8]}};
      2'd2: data__h56748 = {2{soc_clint_s_xactor_f_wr_data_D_OUT[39:8]}};
      2'd3: data__h56748 = soc_clint_s_xactor_f_wr_data_D_OUT[71:8];
    endcase
  end
  always@(soc_clint_s_xactor_f_wr_addr_D_OUT)
  begin
    case (soc_clint_s_xactor_f_wr_addr_D_OUT[1:0])
      2'd0: mask__h56747 = 64'h00000000000000FF;
      2'd1: mask__h56747 = 64'h000000000000FFFF;
      2'd2: mask__h56747 = 64'h00000000FFFFFFFF;
      2'd3: mask__h56747 = 64'hFFFFFFFFFFFFFFFF;
    endcase
  end
  always@(soc_clint_s_xactor_f_rd_addr_D_OUT or
	  temp__h46605 or temp___1__h47250 or temp__h46821 or temp__h56130)
  begin
    case (soc_clint_s_xactor_f_rd_addr_D_OUT[1:0])
      2'd0:
	  IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078 =
	      temp___1__h47250;
      2'd1:
	  IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078 =
	      temp__h46821;
      2'd2:
	  IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078 =
	      temp__h56130;
      2'd3:
	  IF_soc_clint_s_xactor_f_rd_addr_first__009_BIT_ETC___d1078 =
	      temp__h46605;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        soc_clint_clint_msip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	soc_clint_clint_mtip <= `BSV_ASSIGNMENT_DELAY 1'd0;
	soc_clint_clint_rg_tick <= `BSV_ASSIGNMENT_DELAY 4'd0;
	soc_clint_clint_rgmtime <= `BSV_ASSIGNMENT_DELAY 64'd0;
	soc_clint_clint_rgmtimecmp <= `BSV_ASSIGNMENT_DELAY 64'd0;
	soc_uart_user_ifc_baud_value <= `BSV_ASSIGNMENT_DELAY 16'd5;
	soc_uart_user_ifc_uart_fifoRecv_countReg <= `BSV_ASSIGNMENT_DELAY
	    5'd0;
	soc_uart_user_ifc_uart_fifoXmit_countReg <= `BSV_ASSIGNMENT_DELAY
	    5'd0;
	soc_uart_user_ifc_uart_rRecvData <= `BSV_ASSIGNMENT_DELAY 1'd1;
      end
    else
      begin
        if (soc_clint_clint_msip_EN)
	  soc_clint_clint_msip <= `BSV_ASSIGNMENT_DELAY
	      soc_clint_clint_msip_D_IN;
	if (soc_clint_clint_mtip_EN)
	  soc_clint_clint_mtip <= `BSV_ASSIGNMENT_DELAY
	      soc_clint_clint_mtip_D_IN;
	if (soc_clint_clint_rg_tick_EN)
	  soc_clint_clint_rg_tick <= `BSV_ASSIGNMENT_DELAY
	      soc_clint_clint_rg_tick_D_IN;
	if (soc_clint_clint_rgmtime_EN)
	  soc_clint_clint_rgmtime <= `BSV_ASSIGNMENT_DELAY
	      soc_clint_clint_rgmtime_D_IN;
	if (soc_clint_clint_rgmtimecmp_EN)
	  soc_clint_clint_rgmtimecmp <= `BSV_ASSIGNMENT_DELAY
	      soc_clint_clint_rgmtimecmp_D_IN;
	if (soc_uart_user_ifc_baud_value_EN)
	  soc_uart_user_ifc_baud_value <= `BSV_ASSIGNMENT_DELAY
	      soc_uart_user_ifc_baud_value_D_IN;
	if (soc_uart_user_ifc_uart_fifoRecv_countReg_EN)
	  soc_uart_user_ifc_uart_fifoRecv_countReg <= `BSV_ASSIGNMENT_DELAY
	      soc_uart_user_ifc_uart_fifoRecv_countReg_D_IN;
	if (soc_uart_user_ifc_uart_fifoXmit_countReg_EN)
	  soc_uart_user_ifc_uart_fifoXmit_countReg <= `BSV_ASSIGNMENT_DELAY
	      soc_uart_user_ifc_uart_fifoXmit_countReg_D_IN;
	if (soc_uart_user_ifc_uart_rRecvData_EN)
	  soc_uart_user_ifc_uart_rRecvData <= `BSV_ASSIGNMENT_DELAY
	      soc_uart_user_ifc_uart_rRecvData_D_IN;
      end
    if (soc_uart_user_ifc_uart_vrRecvBuffer_0_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_0 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_0_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_1_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_1 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_1_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_2_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_2 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_2_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_3_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_3 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_3_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_4_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_4 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_4_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_5_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_5 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_5_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_6_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_6 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_6_D_IN;
    if (soc_uart_user_ifc_uart_vrRecvBuffer_7_EN)
      soc_uart_user_ifc_uart_vrRecvBuffer_7 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrRecvBuffer_7_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_0_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_0 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_0_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_1_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_1 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_1_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_2_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_2 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_2_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_3_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_3 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_3_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_4_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_4 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_4_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_5_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_5 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_5_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_6_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_6 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_6_D_IN;
    if (soc_uart_user_ifc_uart_vrXmitBuffer_7_EN)
      soc_uart_user_ifc_uart_vrXmitBuffer_7 <= `BSV_ASSIGNMENT_DELAY
	  soc_uart_user_ifc_uart_vrXmitBuffer_7_D_IN;
  end

  always@(posedge CLK or `BSV_RESET_EDGE RST_N)
  if (RST_N == `BSV_RESET_VALUE)
    begin
      soc_uart_user_ifc_uart_rRecvBitCount <= `BSV_ASSIGNMENT_DELAY 4'd0;
      soc_uart_user_ifc_uart_rRecvCellCount <= `BSV_ASSIGNMENT_DELAY 4'd0;
      soc_uart_user_ifc_uart_rRecvParity <= `BSV_ASSIGNMENT_DELAY 1'd0;
      soc_uart_user_ifc_uart_rRecvState <= `BSV_ASSIGNMENT_DELAY 3'd0;
      soc_uart_user_ifc_uart_rXmitBitCount <= `BSV_ASSIGNMENT_DELAY 4'd0;
      soc_uart_user_ifc_uart_rXmitCellCount <= `BSV_ASSIGNMENT_DELAY 4'd0;
      soc_uart_user_ifc_uart_rXmitDataOut <= `BSV_ASSIGNMENT_DELAY 1'd1;
      soc_uart_user_ifc_uart_rXmitParity <= `BSV_ASSIGNMENT_DELAY 1'd0;
      soc_uart_user_ifc_uart_rXmitState <= `BSV_ASSIGNMENT_DELAY 3'd0;
    end
  else
    begin
      if (soc_uart_user_ifc_uart_rRecvBitCount_EN)
	soc_uart_user_ifc_uart_rRecvBitCount <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rRecvBitCount_D_IN;
      if (soc_uart_user_ifc_uart_rRecvCellCount_EN)
	soc_uart_user_ifc_uart_rRecvCellCount <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rRecvCellCount_D_IN;
      if (soc_uart_user_ifc_uart_rRecvParity_EN)
	soc_uart_user_ifc_uart_rRecvParity <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rRecvParity_D_IN;
      if (soc_uart_user_ifc_uart_rRecvState_EN)
	soc_uart_user_ifc_uart_rRecvState <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rRecvState_D_IN;
      if (soc_uart_user_ifc_uart_rXmitBitCount_EN)
	soc_uart_user_ifc_uart_rXmitBitCount <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rXmitBitCount_D_IN;
      if (soc_uart_user_ifc_uart_rXmitCellCount_EN)
	soc_uart_user_ifc_uart_rXmitCellCount <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rXmitCellCount_D_IN;
      if (soc_uart_user_ifc_uart_rXmitDataOut_EN)
	soc_uart_user_ifc_uart_rXmitDataOut <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rXmitDataOut_D_IN;
      if (soc_uart_user_ifc_uart_rXmitParity_EN)
	soc_uart_user_ifc_uart_rXmitParity <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rXmitParity_D_IN;
      if (soc_uart_user_ifc_uart_rXmitState_EN)
	soc_uart_user_ifc_uart_rXmitState <= `BSV_ASSIGNMENT_DELAY
	    soc_uart_user_ifc_uart_rXmitState_D_IN;
    end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    soc_clint_clint_msip = 1'h0;
    soc_clint_clint_mtip = 1'h0;
    soc_clint_clint_rg_tick = 4'hA;
    soc_clint_clint_rgmtime = 64'hAAAAAAAAAAAAAAAA;
    soc_clint_clint_rgmtimecmp = 64'hAAAAAAAAAAAAAAAA;
    soc_uart_user_ifc_baud_value = 16'hAAAA;
    soc_uart_user_ifc_uart_fifoRecv_countReg = 5'h0A;
    soc_uart_user_ifc_uart_fifoXmit_countReg = 5'h0A;
    soc_uart_user_ifc_uart_rRecvBitCount = 4'hA;
    soc_uart_user_ifc_uart_rRecvCellCount = 4'hA;
    soc_uart_user_ifc_uart_rRecvData = 1'h0;
    soc_uart_user_ifc_uart_rRecvParity = 1'h0;
    soc_uart_user_ifc_uart_rRecvState = 3'h2;
    soc_uart_user_ifc_uart_rXmitBitCount = 4'hA;
    soc_uart_user_ifc_uart_rXmitCellCount = 4'hA;
    soc_uart_user_ifc_uart_rXmitDataOut = 1'h0;
    soc_uart_user_ifc_uart_rXmitParity = 1'h0;
    soc_uart_user_ifc_uart_rXmitState = 3'h2;
    soc_uart_user_ifc_uart_vrRecvBuffer_0 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_1 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_2 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_3 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_4 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_5 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_6 = 1'h0;
    soc_uart_user_ifc_uart_vrRecvBuffer_7 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_0 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_1 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_2 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_3 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_4 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_5 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_6 = 1'h0;
    soc_uart_user_ifc_uart_vrXmitBuffer_7 = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule  // mkFormalWrapper

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:12 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// get_inputs                     O   138
// RDY_get_inputs                 O     1 const
// delayed_output                 O   138
// RDY_delayed_output             O     1
// CLK                            I     1 clock
// RST_N                          I     1 reset
// get_inputs_operand1            I    64
// get_inputs_operand2            I    64
// get_inputs_funct3              I     3
// get_inputs_word32              I     1
// EN_get_inputs                  I     1
// EN_delayed_output              I     1 unused
//
// Combinational paths from inputs to outputs:
//   (get_inputs_operand1,
//    get_inputs_operand2,
//    get_inputs_funct3,
//    get_inputs_word32) -> get_inputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkmuldiv(CLK,
		RST_N,

		get_inputs_operand1,
		get_inputs_operand2,
		get_inputs_funct3,
		get_inputs_word32,
		EN_get_inputs,
		get_inputs,
		RDY_get_inputs,

		EN_delayed_output,
		delayed_output,
		RDY_delayed_output);
  input  CLK;
  input  RST_N;

  // actionvalue method get_inputs
  input  [63 : 0] get_inputs_operand1;
  input  [63 : 0] get_inputs_operand2;
  input  [2 : 0] get_inputs_funct3;
  input  get_inputs_word32;
  input  EN_get_inputs;
  output [137 : 0] get_inputs;
  output RDY_get_inputs;

  // actionvalue method delayed_output
  input  EN_delayed_output;
  output [137 : 0] delayed_output;
  output RDY_delayed_output;

  // signals for module outputs
  wire [137 : 0] delayed_output, get_inputs;
  wire RDY_delayed_output, RDY_get_inputs;

  // register mul_div
  reg mul_div;
  wire mul_div_D_IN, mul_div_EN;

  // register mult_reg_a
  reg [127 : 0] mult_reg_a;
  wire [127 : 0] mult_reg_a_D_IN;
  wire mult_reg_a_EN;

  // register mult_reg_b
  reg [127 : 0] mult_reg_b;
  wire [127 : 0] mult_reg_b_D_IN;
  wire mult_reg_b_EN;

  // register rg_complement
  reg rg_complement;
  reg rg_complement_D_IN;
  wire rg_complement_EN;

  // register rg_count
  reg [6 : 0] rg_count;
  wire [6 : 0] rg_count_D_IN;
  wire rg_count_EN;

  // register rg_sign_op1
  reg rg_sign_op1;
  wire rg_sign_op1_D_IN, rg_sign_op1_EN;

  // register rg_upperbits
  reg rg_upperbits;
  wire rg_upperbits_D_IN, rg_upperbits_EN;

  // register rg_word32
  reg rg_word32;
  wire rg_word32_D_IN, rg_word32_EN;

  // ports of submodule divider
  wire [63 : 0] divider_get_inputs_op1,
		divider_get_inputs_op2,
		divider_quo_rem;
  wire divider_EN_get_inputs, divider_get_inputs_qr;

  // rule scheduling signals
  wire CAN_FIRE_RL_increment_counter,
       CAN_FIRE_delayed_output,
       CAN_FIRE_get_inputs,
       WILL_FIRE_RL_increment_counter,
       WILL_FIRE_delayed_output,
       WILL_FIRE_get_inputs;

  // inputs to muxes for submodule ports
  wire [6 : 0] MUX_rg_count_write_1__VAL_2;
  wire MUX_rg_count_write_1__SEL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d102;
  reg TASK_testplusargs___d103;
  reg TASK_testplusargs___d104;
  reg [63 : 0] v__h2313;
  reg TASK_testplusargs___d72;
  reg TASK_testplusargs___d73;
  reg TASK_testplusargs___d74;
  reg [63 : 0] v__h1086;
  reg TASK_testplusargs___d13;
  reg TASK_testplusargs___d14;
  reg TASK_testplusargs___d15;
  reg [63 : 0] v__h482;
  reg TASK_testplusargs___d25;
  reg TASK_testplusargs___d26;
  reg TASK_testplusargs___d27;
  reg [63 : 0] v__h630;
  reg rg_count_EQ_8_AND_NOT_mul_div_OR_rg_count_EQ_6_ETC___d18;
  reg NOT_rg_count_EQ_8_0_OR_mul_div_1_AND_NOT_rg_co_ETC___d30;
  reg NOT_get_inputs_funct3_BIT_2_2_8_AND_TASK_testp_ETC___d77;
  // synopsys translate_on

  // remaining internal signals
  wire [255 : 0] mult_reg_a_26_MUL_mult_reg_b_27___d128;
  wire [127 : 0] _theResult____h2244, reslt___1__h2432, reslt__h2243;
  wire [63 : 0] IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38,
		IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44,
		_theResult_____3_fst__h1845,
		_theResult___fst__h897,
		_theResult___snd__h898,
		default_out___1__h2158,
		default_out__h1785,
		op1__h850,
		op2__h851,
		product__h2245,
		t1__h848,
		t2__h849,
		x__h2154,
		y_avValue_fst__h1777;
  wire [31 : 0] default_out785_BITS_31_TO_0__q3,
		get_inputs_operand1_BITS_31_TO_0__q1,
		get_inputs_operand2_BITS_31_TO_0__q2,
		theResult__244_BITS_31_TO_0__q4;
  wire [6 : 0] x__h724;
  wire IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d88,
       mul_div_AND_rg_upperbits_09_10_AND_rg_compleme_ETC___d118,
       x__h1134,
       x__h1337;

  // actionvalue method get_inputs
  assign get_inputs =
	     { get_inputs_funct3[2] &&
	       IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 ==
	       64'd0,
	       2'd2,
	       x__h2154,
	       64'hAAAAAAAAAAAAAAAA /* unspecified value */ ,
	       6'b101010 /* unspecified value */ ,
	       1'd0 } ;
  assign RDY_get_inputs = 1'd1 ;
  assign CAN_FIRE_get_inputs = 1'd1 ;
  assign WILL_FIRE_get_inputs = EN_get_inputs ;

  // actionvalue method delayed_output
  assign delayed_output =
	     { 3'd6,
	       product__h2245,
	       64'hAAAAAAAAAAAAAAAA /* unspecified value */ ,
	       6'b101010 /* unspecified value */ ,
	       1'd0 } ;
  assign RDY_delayed_output =
	     rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div ;
  assign CAN_FIRE_delayed_output =
	     rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div ;
  assign WILL_FIRE_delayed_output = EN_delayed_output ;

  // submodule divider
  mkrestoring_div divider(.CLK(CLK),
			  .RST_N(RST_N),
			  .get_inputs_op1(divider_get_inputs_op1),
			  .get_inputs_op2(divider_get_inputs_op2),
			  .get_inputs_qr(divider_get_inputs_qr),
			  .EN_get_inputs(divider_EN_get_inputs),
			  .RDY_get_inputs(),
			  .quo_rem(divider_quo_rem),
			  .RDY_quo_rem());

  // rule RL_increment_counter
  assign CAN_FIRE_RL_increment_counter = rg_count != 7'd0 ;
  assign WILL_FIRE_RL_increment_counter =
	     CAN_FIRE_RL_increment_counter && !EN_get_inputs ;

  // inputs to muxes for submodule ports
  assign MUX_rg_count_write_1__SEL_1 =
	     EN_get_inputs &&
	     (!get_inputs_funct3[2] ||
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 !=
	      64'd0) ;
  assign MUX_rg_count_write_1__VAL_2 =
	     (rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div) ?
	       7'd0 :
	       x__h724 ;

  // register mul_div
  assign mul_div_D_IN = get_inputs_funct3[2] ;
  assign mul_div_EN = EN_get_inputs ;

  // register mult_reg_a
  assign mult_reg_a_D_IN = { 64'd0, op1__h850 } ;
  assign mult_reg_a_EN = EN_get_inputs && !get_inputs_funct3[2] ;

  // register mult_reg_b
  assign mult_reg_b_D_IN = { 64'd0, op2__h851 } ;
  assign mult_reg_b_EN = EN_get_inputs && !get_inputs_funct3[2] ;

  // register rg_complement
  always@(get_inputs_funct3 or
	  IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d88 or
	  IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38)
  begin
    case (get_inputs_funct3)
      3'd1, 3'd4:
	  rg_complement_D_IN =
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d88;
      3'd2:
	  rg_complement_D_IN =
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38[63];
      default: rg_complement_D_IN = get_inputs_funct3 == 3'd6;
    endcase
  end
  assign rg_complement_EN = MUX_rg_count_write_1__SEL_1 ;

  // register rg_count
  assign rg_count_D_IN =
	     MUX_rg_count_write_1__SEL_1 ?
	       7'd1 :
	       MUX_rg_count_write_1__VAL_2 ;
  assign rg_count_EN =
	     EN_get_inputs &&
	     (!get_inputs_funct3[2] ||
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 !=
	      64'd0) ||
	     WILL_FIRE_RL_increment_counter ;

  // register rg_sign_op1
  assign rg_sign_op1_D_IN =
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38[63] ;
  assign rg_sign_op1_EN = EN_get_inputs ;

  // register rg_upperbits
  assign rg_upperbits_D_IN =
	     get_inputs_funct3[2] ?
	       get_inputs_funct3[1] :
	       get_inputs_funct3[1:0] != 2'd0 ;
  assign rg_upperbits_EN = MUX_rg_count_write_1__SEL_1 ;

  // register rg_word32
  assign rg_word32_D_IN = get_inputs_word32 ;
  assign rg_word32_EN = MUX_rg_count_write_1__SEL_1 ;

  // submodule divider
  assign divider_get_inputs_op1 = op1__h850 ;
  assign divider_get_inputs_op2 = op2__h851 ;
  assign divider_get_inputs_qr = get_inputs_funct3[1] ;
  assign divider_EN_get_inputs =
	     EN_get_inputs && get_inputs_funct3[2] &&
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 !=
	     64'd0 ;

  // remaining internal signals
  assign IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38 =
	     get_inputs_word32 ?
	       _theResult___fst__h897 :
	       get_inputs_operand1 ;
  assign IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 =
	     get_inputs_word32 ?
	       _theResult___snd__h898 :
	       get_inputs_operand2 ;
  assign IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d88 =
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38[63] ^
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44[63] ;
  assign _theResult_____3_fst__h1845 =
	     get_inputs_funct3[1] ?
	       IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38 :
	       64'hFFFFFFFFFFFFFFFF ;
  assign _theResult____h2244 =
	     (mul_div_AND_rg_upperbits_09_10_AND_rg_compleme_ETC___d118 ||
	      mul_div && rg_complement && !rg_upperbits ||
	      !mul_div && rg_complement) ?
	       reslt___1__h2432 :
	       reslt__h2243 ;
  assign _theResult___fst__h897 =
	     get_inputs_funct3[0] ?
	       { 32'd0, get_inputs_operand1[31:0] } :
	       { {32{get_inputs_operand1_BITS_31_TO_0__q1[31]}},
		 get_inputs_operand1_BITS_31_TO_0__q1 } ;
  assign _theResult___snd__h898 =
	     get_inputs_funct3[0] ?
	       { 32'd0, get_inputs_operand2[31:0] } :
	       { {32{get_inputs_operand2_BITS_31_TO_0__q2[31]}},
		 get_inputs_operand2_BITS_31_TO_0__q2 } ;
  assign default_out785_BITS_31_TO_0__q3 = default_out__h1785[31:0] ;
  assign default_out___1__h2158 =
	     { {32{default_out785_BITS_31_TO_0__q3[31]}},
	       default_out785_BITS_31_TO_0__q3 } ;
  assign default_out__h1785 =
	     get_inputs_funct3[2] ?
	       y_avValue_fst__h1777 :
	       64'hFFFFFFFFFFFFFFFF ;
  assign get_inputs_operand1_BITS_31_TO_0__q1 = get_inputs_operand1[31:0] ;
  assign get_inputs_operand2_BITS_31_TO_0__q2 = get_inputs_operand2[31:0] ;
  assign mul_div_AND_rg_upperbits_09_10_AND_rg_compleme_ETC___d118 =
	     mul_div && rg_upperbits && rg_complement &&
	     divider_quo_rem[63] != rg_sign_op1 ;
  assign mult_reg_a_26_MUL_mult_reg_b_27___d128 = mult_reg_a * mult_reg_b ;
  assign op1__h850 =
	     (t1__h848 ^
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38) +
	     { 63'd0, x__h1134 } ;
  assign op2__h851 =
	     (t2__h849 ^
	      IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44) +
	     { 63'd0, x__h1337 } ;
  assign product__h2245 =
	     rg_word32 ?
	       { {32{theResult__244_BITS_31_TO_0__q4[31]}},
		 theResult__244_BITS_31_TO_0__q4 } :
	       ((!mul_div && rg_upperbits) ?
		  _theResult____h2244[127:64] :
		  _theResult____h2244[63:0]) ;
  assign reslt___1__h2432 = ~reslt__h2243 + 128'd1 ;
  assign reslt__h2243 =
	     mul_div ?
	       { 64'd0, divider_quo_rem } :
	       mult_reg_a_26_MUL_mult_reg_b_27___d128[127:0] ;
  assign t1__h848 = {64{x__h1134}} ;
  assign t2__h849 = {64{x__h1337}} ;
  assign theResult__244_BITS_31_TO_0__q4 = _theResult____h2244[31:0] ;
  assign x__h1134 =
	     !get_inputs_funct3[2] &&
	     get_inputs_funct3[0] ^ get_inputs_funct3[1] &&
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38[63] ||
	     get_inputs_funct3[2] && !get_inputs_funct3[0] &&
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d38[63] ;
  assign x__h1337 =
	     !get_inputs_funct3[2] && get_inputs_funct3[1:0] == 2'd1 &&
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44[63] ||
	     get_inputs_funct3[2] && !get_inputs_funct3[0] &&
	     IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44[63] ;
  assign x__h2154 =
	     get_inputs_word32 ? default_out___1__h2158 : default_out__h1785 ;
  assign x__h724 = rg_count + 7'd1 ;
  assign y_avValue_fst__h1777 =
	     (IF_get_inputs_word32_THEN_IF_get_inputs_funct3_ETC___d44 ==
	      64'd0) ?
	       _theResult_____3_fst__h1845 :
	       64'hFFFFFFFFFFFFFFFF ;

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        mul_div <= `BSV_ASSIGNMENT_DELAY 1'd0;
	mult_reg_a <= `BSV_ASSIGNMENT_DELAY 128'd0;
	mult_reg_b <= `BSV_ASSIGNMENT_DELAY 128'd0;
	rg_complement <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_count <= `BSV_ASSIGNMENT_DELAY 7'd0;
	rg_sign_op1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_upperbits <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_word32 <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (mul_div_EN) mul_div <= `BSV_ASSIGNMENT_DELAY mul_div_D_IN;
	if (mult_reg_a_EN)
	  mult_reg_a <= `BSV_ASSIGNMENT_DELAY mult_reg_a_D_IN;
	if (mult_reg_b_EN)
	  mult_reg_b <= `BSV_ASSIGNMENT_DELAY mult_reg_b_D_IN;
	if (rg_complement_EN)
	  rg_complement <= `BSV_ASSIGNMENT_DELAY rg_complement_D_IN;
	if (rg_count_EN) rg_count <= `BSV_ASSIGNMENT_DELAY rg_count_D_IN;
	if (rg_sign_op1_EN)
	  rg_sign_op1 <= `BSV_ASSIGNMENT_DELAY rg_sign_op1_D_IN;
	if (rg_upperbits_EN)
	  rg_upperbits <= `BSV_ASSIGNMENT_DELAY rg_upperbits_D_IN;
	if (rg_word32_EN) rg_word32 <= `BSV_ASSIGNMENT_DELAY rg_word32_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    mul_div = 1'h0;
    mult_reg_a = 128'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    mult_reg_b = 128'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    rg_complement = 1'h0;
    rg_count = 7'h2A;
    rg_sign_op1 = 1'h0;
    rg_upperbits = 1'h0;
    rg_word32 = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output)
	begin
	  TASK_testplusargs___d102 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output)
	begin
	  TASK_testplusargs___d103 = $test$plusargs("mmuldiv");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output)
	begin
	  TASK_testplusargs___d104 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output)
	begin
	  v__h2313 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output &&
	  (TASK_testplusargs___d102 ||
	   TASK_testplusargs___d103 && TASK_testplusargs___d104))
	$write("[%10d", v__h2313, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output &&
	  (TASK_testplusargs___d102 ||
	   TASK_testplusargs___d103 && TASK_testplusargs___d104))
	$write("MULDIV: Responding with DelayedOut: %h", product__h2245);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_delayed_output &&
	  (TASK_testplusargs___d102 ||
	   TASK_testplusargs___d103 && TASK_testplusargs___d104))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs && !get_inputs_funct3[2])
	begin
	  TASK_testplusargs___d72 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs && !get_inputs_funct3[2])
	begin
	  TASK_testplusargs___d73 = $test$plusargs("mmuldiv");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs && !get_inputs_funct3[2])
	begin
	  TASK_testplusargs___d74 = $test$plusargs("l0");
	  #0;
	end
    NOT_get_inputs_funct3_BIT_2_2_8_AND_TASK_testp_ETC___d77 =
	!get_inputs_funct3[2] &&
	(TASK_testplusargs___d72 ||
	 TASK_testplusargs___d73 && TASK_testplusargs___d74);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs && !get_inputs_funct3[2])
	begin
	  v__h1086 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs &&
	  NOT_get_inputs_funct3_BIT_2_2_8_AND_TASK_testp_ETC___d77)
	$write("[%10d", v__h1086, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs &&
	  NOT_get_inputs_funct3_BIT_2_2_8_AND_TASK_testp_ETC___d77)
	$write("MULDIV : Inps to Mul. A:%h B:%h f3: %b",
	       op1__h850,
	       op2__h851,
	       get_inputs_funct3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_get_inputs &&
	  NOT_get_inputs_funct3_BIT_2_2_8_AND_TASK_testp_ETC___d77)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  (rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div))
	begin
	  TASK_testplusargs___d13 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  (rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div))
	begin
	  TASK_testplusargs___d14 = $test$plusargs("mmuldiv");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  (rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div))
	begin
	  TASK_testplusargs___d15 = $test$plusargs("l0");
	  #0;
	end
    rg_count_EQ_8_AND_NOT_mul_div_OR_rg_count_EQ_6_ETC___d18 =
	(rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div) &&
	(TASK_testplusargs___d13 ||
	 TASK_testplusargs___d14 && TASK_testplusargs___d15);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  (rg_count == 7'd8 && !mul_div || rg_count == 7'd65 && mul_div))
	begin
	  v__h482 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  rg_count_EQ_8_AND_NOT_mul_div_OR_rg_count_EQ_6_ETC___d18)
	$write("[%10d", v__h482, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  rg_count_EQ_8_AND_NOT_mul_div_OR_rg_count_EQ_6_ETC___d18)
	$write("MULDIV : got output from Mul/Div. mul_div: %b", mul_div);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  rg_count_EQ_8_AND_NOT_mul_div_OR_rg_count_EQ_6_ETC___d18)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter && (rg_count != 7'd8 || mul_div) &&
	  (rg_count != 7'd65 || !mul_div))
	begin
	  TASK_testplusargs___d25 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter && (rg_count != 7'd8 || mul_div) &&
	  (rg_count != 7'd65 || !mul_div))
	begin
	  TASK_testplusargs___d26 = $test$plusargs("mmuldiv");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter && (rg_count != 7'd8 || mul_div) &&
	  (rg_count != 7'd65 || !mul_div))
	begin
	  TASK_testplusargs___d27 = $test$plusargs("l0");
	  #0;
	end
    NOT_rg_count_EQ_8_0_OR_mul_div_1_AND_NOT_rg_co_ETC___d30 =
	(rg_count != 7'd8 || mul_div) && (rg_count != 7'd65 || !mul_div) &&
	(TASK_testplusargs___d25 ||
	 TASK_testplusargs___d26 && TASK_testplusargs___d27);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter && (rg_count != 7'd8 || mul_div) &&
	  (rg_count != 7'd65 || !mul_div))
	begin
	  v__h630 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  NOT_rg_count_EQ_8_0_OR_mul_div_1_AND_NOT_rg_co_ETC___d30)
	$write("[%10d", v__h630, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  NOT_rg_count_EQ_8_0_OR_mul_div_1_AND_NOT_rg_co_ETC___d30)
	$write("MULDIV : Waiting for mul/div to respond. Count: %d",
	       rg_count);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_increment_counter &&
	  NOT_rg_count_EQ_8_0_OR_mul_div_1_AND_NOT_rg_co_ETC___d30)
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkmuldiv

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:12 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// RDY_get_inputs                 O     1 const
// quo_rem                        O    64
// RDY_quo_rem                    O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// get_inputs_op1                 I    64
// get_inputs_op2                 I    64 reg
// get_inputs_qr                  I     1 reg
// EN_get_inputs                  I     1
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkrestoring_div(CLK,
		       RST_N,

		       get_inputs_op1,
		       get_inputs_op2,
		       get_inputs_qr,
		       EN_get_inputs,
		       RDY_get_inputs,

		       quo_rem,
		       RDY_quo_rem);
  input  CLK;
  input  RST_N;

  // action method get_inputs
  input  [63 : 0] get_inputs_op1;
  input  [63 : 0] get_inputs_op2;
  input  get_inputs_qr;
  input  EN_get_inputs;
  output RDY_get_inputs;

  // value method quo_rem
  output [63 : 0] quo_rem;
  output RDY_quo_rem;

  // signals for module outputs
  wire [63 : 0] quo_rem;
  wire RDY_get_inputs, RDY_quo_rem;

  // register partial
  reg [128 : 0] partial;
  wire [128 : 0] partial_D_IN;
  wire partial_EN;

  // register quotient_remainder
  reg quotient_remainder;
  wire quotient_remainder_D_IN, quotient_remainder_EN;

  // register rg_op2
  reg [63 : 0] rg_op2;
  wire [63 : 0] rg_op2_D_IN;
  wire rg_op2_EN;

  // rule scheduling signals
  wire CAN_FIRE_RL_single_step_div,
       CAN_FIRE_get_inputs,
       WILL_FIRE_RL_single_step_div,
       WILL_FIRE_get_inputs;

  // inputs to muxes for submodule ports
  wire [128 : 0] MUX_partial_write_1__VAL_1, MUX_partial_write_1__VAL_2;

  // remaining internal signals
  wire [128 : 0] x__h322;
  wire [63 : 0] x_BITS_63_TO_0___h323;

  // action method get_inputs
  assign RDY_get_inputs = 1'd1 ;
  assign CAN_FIRE_get_inputs = 1'd1 ;
  assign WILL_FIRE_get_inputs = EN_get_inputs ;

  // value method quo_rem
  assign quo_rem = quotient_remainder ? partial[127:64] : partial[63:0] ;
  assign RDY_quo_rem = 1'd1 ;

  // rule RL_single_step_div
  assign CAN_FIRE_RL_single_step_div = 1'd1 ;
  assign WILL_FIRE_RL_single_step_div = 1'd1 ;

  // inputs to muxes for submodule ports
  assign MUX_partial_write_1__VAL_1 = { 65'd0, get_inputs_op1 } ;
  module_singlestep instance_singlestep_0(.singlestep_remainder(x__h322[128:64]),
					  .singlestep_quotient(x_BITS_63_TO_0___h323),
					  .singlestep_divisor(rg_op2),
					  .singlestep(MUX_partial_write_1__VAL_2));

  // register partial
  assign partial_D_IN =
	     EN_get_inputs ?
	       MUX_partial_write_1__VAL_1 :
	       MUX_partial_write_1__VAL_2 ;
  assign partial_EN = 1'b1 ;

  // register quotient_remainder
  assign quotient_remainder_D_IN = get_inputs_qr ;
  assign quotient_remainder_EN = EN_get_inputs ;

  // register rg_op2
  assign rg_op2_D_IN = get_inputs_op2 ;
  assign rg_op2_EN = EN_get_inputs ;

  // remaining internal signals
  assign x_BITS_63_TO_0___h323 = partial[63:0] ;
  assign x__h322 = partial ;

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        partial <= `BSV_ASSIGNMENT_DELAY 129'd0;
	quotient_remainder <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_op2 <= `BSV_ASSIGNMENT_DELAY 64'd0;
      end
    else
      begin
        if (partial_EN) partial <= `BSV_ASSIGNMENT_DELAY partial_D_IN;
	if (quotient_remainder_EN)
	  quotient_remainder <= `BSV_ASSIGNMENT_DELAY quotient_remainder_D_IN;
	if (rg_op2_EN) rg_op2 <= `BSV_ASSIGNMENT_DELAY rg_op2_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    partial = 129'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    quotient_remainder = 1'h0;
    rg_op2 = 64'hAAAAAAAAAAAAAAAA;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule  // mkrestoring_div

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:16 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// inst_request_get               O    66
// RDY_inst_request_get           O     1
// RDY_inst_response_put          O     1 reg
// memory_request_get             O   139
// RDY_memory_request_get         O     1 reg
// RDY_memory_response_put        O     1 const
// RDY_clint_msip                 O     1 const
// RDY_clint_mtip                 O     1 const
// RDY_clint_mtime                O     1 const
// RDY_ext_interrupt              O     1 const
// dump_get                       O   167
// RDY_dump_get                   O     1 reg
// mv_curr_priv                   O     2
// RDY_mv_curr_priv               O     1 const
// mv_trap                        O     1
// RDY_mv_trap                    O     1 const
// mv_pmp_cfg                     O    32 reg
// RDY_mv_pmp_cfg                 O     1 const
// mv_pmp_addr                    O   120 reg
// RDY_mv_pmp_addr                O     1 const
// resetpc                        I    64
// CLK                            I     1 clock
// RST_N                          I     1 reset
// inst_response_put              I    35 reg
// memory_response_put            I    66
// clint_msip_intrpt              I     1 reg
// clint_mtip_intrpt              I     1 reg
// clint_mtime_c_mtime            I    64 reg
// ext_interrupt_intrpt           I     1 reg
// EN_inst_response_put           I     1
// EN_memory_response_put         I     1
// EN_clint_msip                  I     1
// EN_clint_mtip                  I     1
// EN_clint_mtime                 I     1
// EN_ext_interrupt               I     1
// EN_inst_request_get            I     1
// EN_memory_request_get          I     1
// EN_dump_get                    I     1
//
// Combinational paths from inputs to outputs:
//   EN_dump_get -> mv_trap
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkriscv(resetpc,
	       CLK,
	       RST_N,

	       EN_inst_request_get,
	       inst_request_get,
	       RDY_inst_request_get,

	       inst_response_put,
	       EN_inst_response_put,
	       RDY_inst_response_put,

	       EN_memory_request_get,
	       memory_request_get,
	       RDY_memory_request_get,

	       memory_response_put,
	       EN_memory_response_put,
	       RDY_memory_response_put,

	       clint_msip_intrpt,
	       EN_clint_msip,
	       RDY_clint_msip,

	       clint_mtip_intrpt,
	       EN_clint_mtip,
	       RDY_clint_mtip,

	       clint_mtime_c_mtime,
	       EN_clint_mtime,
	       RDY_clint_mtime,

	       ext_interrupt_intrpt,
	       EN_ext_interrupt,
	       RDY_ext_interrupt,

	       EN_dump_get,
	       dump_get,
	       RDY_dump_get,

	       mv_curr_priv,
	       RDY_mv_curr_priv,

	       mv_trap,
	       RDY_mv_trap,

	       mv_pmp_cfg,
	       RDY_mv_pmp_cfg,

	       mv_pmp_addr,
	       RDY_mv_pmp_addr);
  input  [63 : 0] resetpc;
  input  CLK;
  input  RST_N;

  // actionvalue method inst_request_get
  input  EN_inst_request_get;
  output [65 : 0] inst_request_get;
  output RDY_inst_request_get;

  // action method inst_response_put
  input  [34 : 0] inst_response_put;
  input  EN_inst_response_put;
  output RDY_inst_response_put;

  // actionvalue method memory_request_get
  input  EN_memory_request_get;
  output [138 : 0] memory_request_get;
  output RDY_memory_request_get;

  // action method memory_response_put
  input  [65 : 0] memory_response_put;
  input  EN_memory_response_put;
  output RDY_memory_response_put;

  // action method clint_msip
  input  clint_msip_intrpt;
  input  EN_clint_msip;
  output RDY_clint_msip;

  // action method clint_mtip
  input  clint_mtip_intrpt;
  input  EN_clint_mtip;
  output RDY_clint_mtip;

  // action method clint_mtime
  input  [63 : 0] clint_mtime_c_mtime;
  input  EN_clint_mtime;
  output RDY_clint_mtime;

  // action method ext_interrupt
  input  ext_interrupt_intrpt;
  input  EN_ext_interrupt;
  output RDY_ext_interrupt;

  // actionvalue method dump_get
  input  EN_dump_get;
  output [166 : 0] dump_get;
  output RDY_dump_get;

  // value method mv_curr_priv
  output [1 : 0] mv_curr_priv;
  output RDY_mv_curr_priv;

  // value method mv_trap
  output mv_trap;
  output RDY_mv_trap;

  // value method mv_pmp_cfg
  output [31 : 0] mv_pmp_cfg;
  output RDY_mv_pmp_cfg;

  // value method mv_pmp_addr
  output [119 : 0] mv_pmp_addr;
  output RDY_mv_pmp_addr;

  // signals for module outputs
  wire [166 : 0] dump_get;
  wire [138 : 0] memory_request_get;
  wire [119 : 0] mv_pmp_addr;
  wire [65 : 0] inst_request_get;
  wire [31 : 0] mv_pmp_cfg;
  wire [1 : 0] mv_curr_priv;
  wire RDY_clint_msip,
       RDY_clint_mtime,
       RDY_clint_mtip,
       RDY_dump_get,
       RDY_ext_interrupt,
       RDY_inst_request_get,
       RDY_inst_response_put,
       RDY_memory_request_get,
       RDY_memory_response_put,
       RDY_mv_curr_priv,
       RDY_mv_pmp_addr,
       RDY_mv_pmp_cfg,
       RDY_mv_trap,
       mv_trap;

  // ports of submodule fifof
  wire [127 : 0] fifof_D_IN, fifof_D_OUT;
  wire fifof_CLR, fifof_DEQ, fifof_EMPTY_N, fifof_ENQ, fifof_FULL_N;

  // ports of submodule fifof_1
  wire [65 : 0] fifof_1_D_IN, fifof_1_D_OUT;
  wire fifof_1_CLR, fifof_1_DEQ, fifof_1_EMPTY_N, fifof_1_ENQ, fifof_1_FULL_N;

  // ports of submodule fifof_2
  wire [64 : 0] fifof_2_D_IN, fifof_2_D_OUT;
  wire fifof_2_CLR, fifof_2_DEQ, fifof_2_EMPTY_N, fifof_2_ENQ, fifof_2_FULL_N;

  // ports of submodule fifof_3
  wire [69 : 0] fifof_3_D_IN, fifof_3_D_OUT;
  wire fifof_3_CLR, fifof_3_DEQ, fifof_3_EMPTY_N, fifof_3_ENQ, fifof_3_FULL_N;

  // ports of submodule fifof_4
  wire [82 : 0] fifof_4_D_IN, fifof_4_D_OUT;
  wire fifof_4_CLR, fifof_4_DEQ, fifof_4_EMPTY_N, fifof_4_ENQ, fifof_4_FULL_N;

  // ports of submodule fifof_5
  wire [95 : 0] fifof_5_D_IN, fifof_5_D_OUT;
  wire fifof_5_CLR, fifof_5_DEQ, fifof_5_EMPTY_N, fifof_5_ENQ, fifof_5_FULL_N;

  // ports of submodule fifof_6
  wire [95 : 0] fifof_6_D_IN, fifof_6_D_OUT;
  wire fifof_6_CLR, fifof_6_DEQ, fifof_6_EMPTY_N, fifof_6_ENQ, fifof_6_FULL_N;

  // ports of submodule stage1
  wire [151 : 0] stage1_ma_csr_decode_c;
  wire [127 : 0] stage1_ma_trigger_data2_t,
		 stage1_tx_stage1_operands_enq_data;
  wire [95 : 0] stage1_tx_stage1_dump_enq_data;
  wire [68 : 0] stage1_commit_rd_put;
  wire [65 : 0] stage1_inst_request_get, stage1_tx_stage1_control_enq_data;
  wire [64 : 0] stage1_tx_stage1_meta_enq_data;
  wire [63 : 0] stage1_ma_flush_newpc;
  wire [43 : 0] stage1_ma_trigger_data1_t;
  wire [34 : 0] stage1_inst_response_put;
  wire [1 : 0] stage1_ma_trigger_enable_t;
  wire stage1_EN_commit_rd_put,
       stage1_EN_inst_request_get,
       stage1_EN_inst_response_put,
       stage1_EN_ma_flush,
       stage1_EN_ma_update_eEpoch,
       stage1_EN_ma_update_wEpoch,
       stage1_RDY_commit_rd_put,
       stage1_RDY_inst_request_get,
       stage1_RDY_inst_response_put,
       stage1_ma_csr_misa_c_c,
       stage1_ma_interrupt_i,
       stage1_tx_stage1_control_enq_ena,
       stage1_tx_stage1_control_enq_rdy_b,
       stage1_tx_stage1_control_notFull_b,
       stage1_tx_stage1_dump_enq_ena,
       stage1_tx_stage1_dump_enq_rdy_b,
       stage1_tx_stage1_dump_notFull_b,
       stage1_tx_stage1_meta_enq_ena,
       stage1_tx_stage1_meta_enq_rdy_b,
       stage1_tx_stage1_meta_notFull_b,
       stage1_tx_stage1_operands_enq_ena,
       stage1_tx_stage1_operands_enq_rdy_b,
       stage1_tx_stage1_operands_notFull_b;

  // ports of submodule stage2
  wire [138 : 0] stage2_memory_request_get;
  wire [127 : 0] stage2_ma_trigger_data2_t, stage2_rx_stage1_operands_first_x;
  wire [95 : 0] stage2_rx_stage1_dump_first_x, stage2_tx_stage3_dump_enq_data;
  wire [82 : 0] stage2_tx_stage3_type_enq_data;
  wire [69 : 0] stage2_operand_fwding_put, stage2_tx_stage3_common_enq_data;
  wire [65 : 0] stage2_rx_stage1_control_first_x;
  wire [64 : 0] stage2_mv_delayed_output, stage2_rx_stage1_meta_first_x;
  wire [63 : 0] stage2_mv_redirection_fst;
  wire [43 : 0] stage2_ma_trigger_data1_t;
  wire [1 : 0] stage2_ma_trigger_enable_t;
  wire stage2_EN_ma_csr_misa_c,
       stage2_EN_ma_update_wEpoch,
       stage2_EN_memory_request_get,
       stage2_EN_operand_fwding_put,
       stage2_RDY_memory_request_get,
       stage2_ma_csr_misa_c_c,
       stage2_mv_redirection_snd,
       stage2_rx_stage1_control_deq_ena,
       stage2_rx_stage1_control_first_deq_rdy_b,
       stage2_rx_stage1_control_notEmpty_b,
       stage2_rx_stage1_dump_deq_ena,
       stage2_rx_stage1_dump_first_deq_rdy_b,
       stage2_rx_stage1_dump_notEmpty_b,
       stage2_rx_stage1_meta_deq_ena,
       stage2_rx_stage1_meta_first_deq_rdy_b,
       stage2_rx_stage1_meta_notEmpty_b,
       stage2_rx_stage1_operands_deq_ena,
       stage2_rx_stage1_operands_first_deq_rdy_b,
       stage2_rx_stage1_operands_notEmpty_b,
       stage2_tx_stage3_common_enq_ena,
       stage2_tx_stage3_common_enq_rdy_b,
       stage2_tx_stage3_common_notFull_b,
       stage2_tx_stage3_dump_enq_ena,
       stage2_tx_stage3_dump_enq_rdy_b,
       stage2_tx_stage3_dump_notFull_b,
       stage2_tx_stage3_type_enq_ena,
       stage2_tx_stage3_type_enq_rdy_b,
       stage2_tx_stage3_type_notFull_b;

  // ports of submodule stage3
  wire [166 : 0] stage3_dump_get;
  wire [151 : 0] stage3_mv_csr_decode;
  wire [127 : 0] stage3_mv_trigger_data2;
  wire [119 : 0] stage3_mv_pmp_addr;
  wire [95 : 0] stage3_rx_stage3_dump_first_x;
  wire [82 : 0] stage3_rx_stage3_type_first_x;
  wire [69 : 0] stage3_operand_fwding_get, stage3_rx_stage3_common_first_x;
  wire [68 : 0] stage3_commit_rd_get;
  wire [65 : 0] stage3_memory_response_put;
  wire [64 : 0] stage3_ma_delayed_output_r;
  wire [63 : 0] stage3_clint_mtime_c_mtime, stage3_flush_fst;
  wire [43 : 0] stage3_mv_trigger_data1;
  wire [31 : 0] stage3_mv_pmp_cfg;
  wire [1 : 0] stage3_mv_curr_priv, stage3_mv_trigger_enable;
  wire stage3_EN_clint_msip,
       stage3_EN_clint_mtime,
       stage3_EN_clint_mtip,
       stage3_EN_commit_rd_get,
       stage3_EN_dump_get,
       stage3_EN_ext_interrupt,
       stage3_EN_ma_delayed_output,
       stage3_EN_memory_response_put,
       stage3_EN_operand_fwding_get,
       stage3_RDY_commit_rd_get,
       stage3_RDY_dump_get,
       stage3_clint_msip_intrpt,
       stage3_clint_mtip_intrpt,
       stage3_ext_interrupt_i,
       stage3_flush_snd,
       stage3_mv_csr_misa_c,
       stage3_mv_interrupt,
       stage3_rx_stage3_common_deq_ena,
       stage3_rx_stage3_common_first_deq_rdy_b,
       stage3_rx_stage3_common_notEmpty_b,
       stage3_rx_stage3_dump_deq_ena,
       stage3_rx_stage3_dump_first_deq_rdy_b,
       stage3_rx_stage3_dump_notEmpty_b,
       stage3_rx_stage3_type_deq_ena,
       stage3_rx_stage3_type_first_deq_rdy_b,
       stage3_rx_stage3_type_notEmpty_b;

  // rule scheduling signals
  wire CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_rdy,
       CAN_FIRE_RL_empty_fifof_to_rxe_connect_ena,
       CAN_FIRE_RL_empty_fifof_to_rxe_connect_first,
       CAN_FIRE_RL_empty_fifof_to_rxe_connect_notEmpty,
       CAN_FIRE_RL_empty_fifof_to_rxe_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_1_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_1_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_2_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_2_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_3_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_3_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_4_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_4_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_5_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_5_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_6_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_6_connect_rdy,
       CAN_FIRE_RL_empty_txe_to_fifof_connect_ena_data,
       CAN_FIRE_RL_empty_txe_to_fifof_connect_notFull,
       CAN_FIRE_RL_empty_txe_to_fifof_connect_rdy,
       CAN_FIRE_RL_flush_from_writeback,
       CAN_FIRE_RL_gen_new_pc,
       CAN_FIRE_RL_mkConnectionGetPut,
       CAN_FIRE_RL_mkConnectionGetPut_1,
       CAN_FIRE_RL_mkConnectionVtoAf,
       CAN_FIRE_RL_mkConnectionVtoAf_1,
       CAN_FIRE_RL_mkConnectionVtoAf_10,
       CAN_FIRE_RL_mkConnectionVtoAf_2,
       CAN_FIRE_RL_mkConnectionVtoAf_3,
       CAN_FIRE_RL_mkConnectionVtoAf_4,
       CAN_FIRE_RL_mkConnectionVtoAf_5,
       CAN_FIRE_RL_mkConnectionVtoAf_6,
       CAN_FIRE_RL_mkConnectionVtoAf_7,
       CAN_FIRE_RL_mkConnectionVtoAf_8,
       CAN_FIRE_RL_mkConnectionVtoAf_9,
       CAN_FIRE_RL_redirection_from_stage2,
       CAN_FIRE_clint_msip,
       CAN_FIRE_clint_mtime,
       CAN_FIRE_clint_mtip,
       CAN_FIRE_dump_get,
       CAN_FIRE_ext_interrupt,
       CAN_FIRE_inst_request_get,
       CAN_FIRE_inst_response_put,
       CAN_FIRE_memory_request_get,
       CAN_FIRE_memory_response_put,
       WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_rdy,
       WILL_FIRE_RL_empty_fifof_to_rxe_connect_ena,
       WILL_FIRE_RL_empty_fifof_to_rxe_connect_first,
       WILL_FIRE_RL_empty_fifof_to_rxe_connect_notEmpty,
       WILL_FIRE_RL_empty_fifof_to_rxe_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_1_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_1_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_2_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_2_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_3_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_3_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_4_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_4_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_5_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_5_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_6_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_6_connect_rdy,
       WILL_FIRE_RL_empty_txe_to_fifof_connect_ena_data,
       WILL_FIRE_RL_empty_txe_to_fifof_connect_notFull,
       WILL_FIRE_RL_empty_txe_to_fifof_connect_rdy,
       WILL_FIRE_RL_flush_from_writeback,
       WILL_FIRE_RL_gen_new_pc,
       WILL_FIRE_RL_mkConnectionGetPut,
       WILL_FIRE_RL_mkConnectionGetPut_1,
       WILL_FIRE_RL_mkConnectionVtoAf,
       WILL_FIRE_RL_mkConnectionVtoAf_1,
       WILL_FIRE_RL_mkConnectionVtoAf_10,
       WILL_FIRE_RL_mkConnectionVtoAf_2,
       WILL_FIRE_RL_mkConnectionVtoAf_3,
       WILL_FIRE_RL_mkConnectionVtoAf_4,
       WILL_FIRE_RL_mkConnectionVtoAf_5,
       WILL_FIRE_RL_mkConnectionVtoAf_6,
       WILL_FIRE_RL_mkConnectionVtoAf_7,
       WILL_FIRE_RL_mkConnectionVtoAf_8,
       WILL_FIRE_RL_mkConnectionVtoAf_9,
       WILL_FIRE_RL_redirection_from_stage2,
       WILL_FIRE_clint_msip,
       WILL_FIRE_clint_mtime,
       WILL_FIRE_clint_mtip,
       WILL_FIRE_dump_get,
       WILL_FIRE_ext_interrupt,
       WILL_FIRE_inst_request_get,
       WILL_FIRE_inst_response_put,
       WILL_FIRE_memory_request_get,
       WILL_FIRE_memory_response_put;

  // remaining internal signals
  reg [21 : 0] CASE_stage3mv_trigger_data1_BITS_21_TO_20_0_s_ETC__q6,
	       CASE_stage3mv_trigger_data1_BITS_43_TO_42_0_s_ETC__q5;
  reg [1 : 0] CASE_IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_fi_ETC__q7,
	      CASE_IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_f_ETC__q8,
	      CASE_stage1tx_stage1_meta_enq_data_BITS_42_TO_ETC__q2,
	      CASE_stage2memory_request_get_BITS_10_TO_9_0__ETC__q1,
	      CASE_stage2tx_stage3_type_enq_data_BITS_67_TO_ETC__q4,
	      CASE_stage2tx_stage3_type_enq_data_BITS_82_TO_ETC__q3,
	      IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57,
	      IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121;

  // actionvalue method inst_request_get
  assign inst_request_get = stage1_inst_request_get ;
  assign RDY_inst_request_get = stage1_RDY_inst_request_get ;
  assign CAN_FIRE_inst_request_get = stage1_RDY_inst_request_get ;
  assign WILL_FIRE_inst_request_get = EN_inst_request_get ;

  // action method inst_response_put
  assign RDY_inst_response_put = stage1_RDY_inst_response_put ;
  assign CAN_FIRE_inst_response_put = stage1_RDY_inst_response_put ;
  assign WILL_FIRE_inst_response_put = EN_inst_response_put ;

  // actionvalue method memory_request_get
  assign memory_request_get =
	     { stage2_memory_request_get[138:11],
	       CASE_stage2memory_request_get_BITS_10_TO_9_0__ETC__q1,
	       stage2_memory_request_get[8:0] } ;
  assign RDY_memory_request_get = stage2_RDY_memory_request_get ;
  assign CAN_FIRE_memory_request_get = stage2_RDY_memory_request_get ;
  assign WILL_FIRE_memory_request_get = EN_memory_request_get ;

  // action method memory_response_put
  assign RDY_memory_response_put = 1'd1 ;
  assign CAN_FIRE_memory_response_put = 1'd1 ;
  assign WILL_FIRE_memory_response_put = EN_memory_response_put ;

  // action method clint_msip
  assign RDY_clint_msip = 1'd1 ;
  assign CAN_FIRE_clint_msip = 1'd1 ;
  assign WILL_FIRE_clint_msip = EN_clint_msip ;

  // action method clint_mtip
  assign RDY_clint_mtip = 1'd1 ;
  assign CAN_FIRE_clint_mtip = 1'd1 ;
  assign WILL_FIRE_clint_mtip = EN_clint_mtip ;

  // action method clint_mtime
  assign RDY_clint_mtime = 1'd1 ;
  assign CAN_FIRE_clint_mtime = 1'd1 ;
  assign WILL_FIRE_clint_mtime = EN_clint_mtime ;

  // action method ext_interrupt
  assign RDY_ext_interrupt = 1'd1 ;
  assign CAN_FIRE_ext_interrupt = 1'd1 ;
  assign WILL_FIRE_ext_interrupt = EN_ext_interrupt ;

  // actionvalue method dump_get
  assign dump_get =
	     { (stage3_dump_get[166:165] == 2'd3) ?
		 stage3_dump_get[166:165] :
		 2'd0,
	       stage3_dump_get[164:0] } ;
  assign RDY_dump_get = stage3_RDY_dump_get ;
  assign CAN_FIRE_dump_get = stage3_RDY_dump_get ;
  assign WILL_FIRE_dump_get = EN_dump_get ;

  // value method mv_curr_priv
  assign mv_curr_priv = stage3_mv_curr_priv ;
  assign RDY_mv_curr_priv = 1'd1 ;

  // value method mv_trap
  assign mv_trap = stage3_flush_snd ;
  assign RDY_mv_trap = 1'd1 ;

  // value method mv_pmp_cfg
  assign mv_pmp_cfg = stage3_mv_pmp_cfg ;
  assign RDY_mv_pmp_cfg = 1'd1 ;

  // value method mv_pmp_addr
  assign mv_pmp_addr = stage3_mv_pmp_addr ;
  assign RDY_mv_pmp_addr = 1'd1 ;

  // submodule fifof
  FIFOL1 #(.width(32'd128)) fifof(.RST(RST_N),
				  .CLK(CLK),
				  .D_IN(fifof_D_IN),
				  .ENQ(fifof_ENQ),
				  .DEQ(fifof_DEQ),
				  .CLR(fifof_CLR),
				  .D_OUT(fifof_D_OUT),
				  .FULL_N(fifof_FULL_N),
				  .EMPTY_N(fifof_EMPTY_N));

  // submodule fifof_1
  FIFOL1 #(.width(32'd66)) fifof_1(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_1_D_IN),
				   .ENQ(fifof_1_ENQ),
				   .DEQ(fifof_1_DEQ),
				   .CLR(fifof_1_CLR),
				   .D_OUT(fifof_1_D_OUT),
				   .FULL_N(fifof_1_FULL_N),
				   .EMPTY_N(fifof_1_EMPTY_N));

  // submodule fifof_2
  FIFOL1 #(.width(32'd65)) fifof_2(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_2_D_IN),
				   .ENQ(fifof_2_ENQ),
				   .DEQ(fifof_2_DEQ),
				   .CLR(fifof_2_CLR),
				   .D_OUT(fifof_2_D_OUT),
				   .FULL_N(fifof_2_FULL_N),
				   .EMPTY_N(fifof_2_EMPTY_N));

  // submodule fifof_3
  FIFOL1 #(.width(32'd70)) fifof_3(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_3_D_IN),
				   .ENQ(fifof_3_ENQ),
				   .DEQ(fifof_3_DEQ),
				   .CLR(fifof_3_CLR),
				   .D_OUT(fifof_3_D_OUT),
				   .FULL_N(fifof_3_FULL_N),
				   .EMPTY_N(fifof_3_EMPTY_N));

  // submodule fifof_4
  FIFOL1 #(.width(32'd83)) fifof_4(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_4_D_IN),
				   .ENQ(fifof_4_ENQ),
				   .DEQ(fifof_4_DEQ),
				   .CLR(fifof_4_CLR),
				   .D_OUT(fifof_4_D_OUT),
				   .FULL_N(fifof_4_FULL_N),
				   .EMPTY_N(fifof_4_EMPTY_N));

  // submodule fifof_5
  FIFOL1 #(.width(32'd96)) fifof_5(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_5_D_IN),
				   .ENQ(fifof_5_ENQ),
				   .DEQ(fifof_5_DEQ),
				   .CLR(fifof_5_CLR),
				   .D_OUT(fifof_5_D_OUT),
				   .FULL_N(fifof_5_FULL_N),
				   .EMPTY_N(fifof_5_EMPTY_N));

  // submodule fifof_6
  FIFOL1 #(.width(32'd96)) fifof_6(.RST(RST_N),
				   .CLK(CLK),
				   .D_IN(fifof_6_D_IN),
				   .ENQ(fifof_6_ENQ),
				   .DEQ(fifof_6_DEQ),
				   .CLR(fifof_6_CLR),
				   .D_OUT(fifof_6_D_OUT),
				   .FULL_N(fifof_6_FULL_N),
				   .EMPTY_N(fifof_6_EMPTY_N));

  // submodule stage1
  mkstage1 stage1(.resetpc(resetpc),
		  .CLK(CLK),
		  .RST_N(RST_N),
		  .commit_rd_put(stage1_commit_rd_put),
		  .inst_response_put(stage1_inst_response_put),
		  .ma_csr_decode_c(stage1_ma_csr_decode_c),
		  .ma_csr_misa_c_c(stage1_ma_csr_misa_c_c),
		  .ma_flush_newpc(stage1_ma_flush_newpc),
		  .ma_interrupt_i(stage1_ma_interrupt_i),
		  .ma_trigger_data1_t(stage1_ma_trigger_data1_t),
		  .ma_trigger_data2_t(stage1_ma_trigger_data2_t),
		  .ma_trigger_enable_t(stage1_ma_trigger_enable_t),
		  .tx_stage1_control_enq_rdy_b(stage1_tx_stage1_control_enq_rdy_b),
		  .tx_stage1_control_notFull_b(stage1_tx_stage1_control_notFull_b),
		  .tx_stage1_dump_enq_rdy_b(stage1_tx_stage1_dump_enq_rdy_b),
		  .tx_stage1_dump_notFull_b(stage1_tx_stage1_dump_notFull_b),
		  .tx_stage1_meta_enq_rdy_b(stage1_tx_stage1_meta_enq_rdy_b),
		  .tx_stage1_meta_notFull_b(stage1_tx_stage1_meta_notFull_b),
		  .tx_stage1_operands_enq_rdy_b(stage1_tx_stage1_operands_enq_rdy_b),
		  .tx_stage1_operands_notFull_b(stage1_tx_stage1_operands_notFull_b),
		  .EN_inst_request_get(stage1_EN_inst_request_get),
		  .EN_inst_response_put(stage1_EN_inst_response_put),
		  .EN_commit_rd_put(stage1_EN_commit_rd_put),
		  .EN_ma_flush(stage1_EN_ma_flush),
		  .EN_ma_update_eEpoch(stage1_EN_ma_update_eEpoch),
		  .EN_ma_update_wEpoch(stage1_EN_ma_update_wEpoch),
		  .inst_request_get(stage1_inst_request_get),
		  .RDY_inst_request_get(stage1_RDY_inst_request_get),
		  .RDY_inst_response_put(stage1_RDY_inst_response_put),
		  .tx_stage1_operands_enq_ena(stage1_tx_stage1_operands_enq_ena),
		  .tx_stage1_operands_enq_data(stage1_tx_stage1_operands_enq_data),
		  .tx_stage1_meta_enq_ena(stage1_tx_stage1_meta_enq_ena),
		  .tx_stage1_meta_enq_data(stage1_tx_stage1_meta_enq_data),
		  .tx_stage1_control_enq_ena(stage1_tx_stage1_control_enq_ena),
		  .tx_stage1_control_enq_data(stage1_tx_stage1_control_enq_data),
		  .tx_stage1_dump_enq_ena(stage1_tx_stage1_dump_enq_ena),
		  .tx_stage1_dump_enq_data(stage1_tx_stage1_dump_enq_data),
		  .RDY_commit_rd_put(stage1_RDY_commit_rd_put),
		  .RDY_ma_update_eEpoch(),
		  .RDY_ma_update_wEpoch());

  // submodule stage2
  mkstage2 stage2(.CLK(CLK),
		  .RST_N(RST_N),
		  .ma_csr_misa_c_c(stage2_ma_csr_misa_c_c),
		  .ma_trigger_data1_t(stage2_ma_trigger_data1_t),
		  .ma_trigger_data2_t(stage2_ma_trigger_data2_t),
		  .ma_trigger_enable_t(stage2_ma_trigger_enable_t),
		  .operand_fwding_put(stage2_operand_fwding_put),
		  .rx_stage1_control_first_deq_rdy_b(stage2_rx_stage1_control_first_deq_rdy_b),
		  .rx_stage1_control_first_x(stage2_rx_stage1_control_first_x),
		  .rx_stage1_control_notEmpty_b(stage2_rx_stage1_control_notEmpty_b),
		  .rx_stage1_dump_first_deq_rdy_b(stage2_rx_stage1_dump_first_deq_rdy_b),
		  .rx_stage1_dump_first_x(stage2_rx_stage1_dump_first_x),
		  .rx_stage1_dump_notEmpty_b(stage2_rx_stage1_dump_notEmpty_b),
		  .rx_stage1_meta_first_deq_rdy_b(stage2_rx_stage1_meta_first_deq_rdy_b),
		  .rx_stage1_meta_first_x(stage2_rx_stage1_meta_first_x),
		  .rx_stage1_meta_notEmpty_b(stage2_rx_stage1_meta_notEmpty_b),
		  .rx_stage1_operands_first_deq_rdy_b(stage2_rx_stage1_operands_first_deq_rdy_b),
		  .rx_stage1_operands_first_x(stage2_rx_stage1_operands_first_x),
		  .rx_stage1_operands_notEmpty_b(stage2_rx_stage1_operands_notEmpty_b),
		  .tx_stage3_common_enq_rdy_b(stage2_tx_stage3_common_enq_rdy_b),
		  .tx_stage3_common_notFull_b(stage2_tx_stage3_common_notFull_b),
		  .tx_stage3_dump_enq_rdy_b(stage2_tx_stage3_dump_enq_rdy_b),
		  .tx_stage3_dump_notFull_b(stage2_tx_stage3_dump_notFull_b),
		  .tx_stage3_type_enq_rdy_b(stage2_tx_stage3_type_enq_rdy_b),
		  .tx_stage3_type_notFull_b(stage2_tx_stage3_type_notFull_b),
		  .EN_memory_request_get(stage2_EN_memory_request_get),
		  .EN_operand_fwding_put(stage2_EN_operand_fwding_put),
		  .EN_ma_update_wEpoch(stage2_EN_ma_update_wEpoch),
		  .EN_ma_csr_misa_c(stage2_EN_ma_csr_misa_c),
		  .rx_stage1_operands_deq_ena(stage2_rx_stage1_operands_deq_ena),
		  .rx_stage1_meta_deq_ena(stage2_rx_stage1_meta_deq_ena),
		  .rx_stage1_control_deq_ena(stage2_rx_stage1_control_deq_ena),
		  .tx_stage3_common_enq_ena(stage2_tx_stage3_common_enq_ena),
		  .tx_stage3_common_enq_data(stage2_tx_stage3_common_enq_data),
		  .tx_stage3_type_enq_ena(stage2_tx_stage3_type_enq_ena),
		  .tx_stage3_type_enq_data(stage2_tx_stage3_type_enq_data),
		  .rx_stage1_dump_deq_ena(stage2_rx_stage1_dump_deq_ena),
		  .tx_stage3_dump_enq_ena(stage2_tx_stage3_dump_enq_ena),
		  .tx_stage3_dump_enq_data(stage2_tx_stage3_dump_enq_data),
		  .memory_request_get(stage2_memory_request_get),
		  .RDY_memory_request_get(stage2_RDY_memory_request_get),
		  .RDY_operand_fwding_put(),
		  .RDY_ma_update_wEpoch(),
		  .RDY_ma_csr_misa_c(),
		  .mv_delayed_output(stage2_mv_delayed_output),
		  .RDY_mv_delayed_output(),
		  .mv_redirection_fst(stage2_mv_redirection_fst),
		  .RDY_mv_redirection_fst(),
		  .mv_redirection_snd(stage2_mv_redirection_snd),
		  .RDY_mv_redirection_snd());

  // submodule stage3
  mkstage3 stage3(.CLK(CLK),
		  .RST_N(RST_N),
		  .clint_msip_intrpt(stage3_clint_msip_intrpt),
		  .clint_mtime_c_mtime(stage3_clint_mtime_c_mtime),
		  .clint_mtip_intrpt(stage3_clint_mtip_intrpt),
		  .ext_interrupt_i(stage3_ext_interrupt_i),
		  .ma_delayed_output_r(stage3_ma_delayed_output_r),
		  .memory_response_put(stage3_memory_response_put),
		  .rx_stage3_common_first_deq_rdy_b(stage3_rx_stage3_common_first_deq_rdy_b),
		  .rx_stage3_common_first_x(stage3_rx_stage3_common_first_x),
		  .rx_stage3_common_notEmpty_b(stage3_rx_stage3_common_notEmpty_b),
		  .rx_stage3_dump_first_deq_rdy_b(stage3_rx_stage3_dump_first_deq_rdy_b),
		  .rx_stage3_dump_first_x(stage3_rx_stage3_dump_first_x),
		  .rx_stage3_dump_notEmpty_b(stage3_rx_stage3_dump_notEmpty_b),
		  .rx_stage3_type_first_deq_rdy_b(stage3_rx_stage3_type_first_deq_rdy_b),
		  .rx_stage3_type_first_x(stage3_rx_stage3_type_first_x),
		  .rx_stage3_type_notEmpty_b(stage3_rx_stage3_type_notEmpty_b),
		  .EN_memory_response_put(stage3_EN_memory_response_put),
		  .EN_commit_rd_get(stage3_EN_commit_rd_get),
		  .EN_operand_fwding_get(stage3_EN_operand_fwding_get),
		  .EN_clint_msip(stage3_EN_clint_msip),
		  .EN_clint_mtip(stage3_EN_clint_mtip),
		  .EN_clint_mtime(stage3_EN_clint_mtime),
		  .EN_ext_interrupt(stage3_EN_ext_interrupt),
		  .EN_dump_get(stage3_EN_dump_get),
		  .EN_ma_delayed_output(stage3_EN_ma_delayed_output),
		  .rx_stage3_common_deq_ena(stage3_rx_stage3_common_deq_ena),
		  .rx_stage3_type_deq_ena(stage3_rx_stage3_type_deq_ena),
		  .rx_stage3_dump_deq_ena(stage3_rx_stage3_dump_deq_ena),
		  .RDY_memory_response_put(),
		  .commit_rd_get(stage3_commit_rd_get),
		  .RDY_commit_rd_get(stage3_RDY_commit_rd_get),
		  .operand_fwding_get(stage3_operand_fwding_get),
		  .RDY_operand_fwding_get(),
		  .flush_fst(stage3_flush_fst),
		  .RDY_flush_fst(),
		  .flush_snd(stage3_flush_snd),
		  .RDY_flush_snd(),
		  .mv_csr_decode(stage3_mv_csr_decode),
		  .RDY_mv_csr_decode(),
		  .mv_csr_misa_c(stage3_mv_csr_misa_c),
		  .RDY_mv_csr_misa_c(),
		  .RDY_clint_msip(),
		  .RDY_clint_mtip(),
		  .RDY_clint_mtime(),
		  .RDY_ext_interrupt(),
		  .csr_updated(),
		  .RDY_csr_updated(),
		  .mv_interrupt(stage3_mv_interrupt),
		  .dump_get(stage3_dump_get),
		  .RDY_dump_get(stage3_RDY_dump_get),
		  .mv_trigger_data1(stage3_mv_trigger_data1),
		  .RDY_mv_trigger_data1(),
		  .mv_trigger_data2(stage3_mv_trigger_data2),
		  .RDY_mv_trigger_data2(),
		  .mv_trigger_enable(stage3_mv_trigger_enable),
		  .RDY_mv_trigger_enable(),
		  .mv_curr_priv(stage3_mv_curr_priv),
		  .RDY_mv_curr_priv(),
		  .RDY_ma_delayed_output(),
		  .mv_pmp_cfg(stage3_mv_pmp_cfg),
		  .RDY_mv_pmp_cfg(),
		  .mv_pmp_addr(stage3_mv_pmp_addr),
		  .RDY_mv_pmp_addr());

  // rule RL_mkConnectionVtoAf
  assign CAN_FIRE_RL_mkConnectionVtoAf = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf = 1'd1 ;

  // rule RL_mkConnectionVtoAf_1
  assign CAN_FIRE_RL_mkConnectionVtoAf_1 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_1 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_2
  assign CAN_FIRE_RL_mkConnectionVtoAf_2 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_2 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_3
  assign CAN_FIRE_RL_mkConnectionVtoAf_3 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_3 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_4
  assign CAN_FIRE_RL_mkConnectionVtoAf_4 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_4 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_5
  assign CAN_FIRE_RL_mkConnectionVtoAf_5 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_5 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_6
  assign CAN_FIRE_RL_mkConnectionVtoAf_6 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_6 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_7
  assign CAN_FIRE_RL_mkConnectionVtoAf_7 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_7 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_8
  assign CAN_FIRE_RL_mkConnectionVtoAf_8 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_8 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_9
  assign CAN_FIRE_RL_mkConnectionVtoAf_9 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_9 = 1'd1 ;

  // rule RL_mkConnectionVtoAf_10
  assign CAN_FIRE_RL_mkConnectionVtoAf_10 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionVtoAf_10 = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_connect_first = fifof_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_connect_first = fifof_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_1_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_1_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_1_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_first = fifof_1_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_first = fifof_1_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_2_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_2_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_2_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_first = fifof_2_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_first = fifof_2_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_3_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_3_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_3_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_first = fifof_3_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_first = fifof_3_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_4_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_4_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_4_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_first = fifof_4_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_first = fifof_4_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_5_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_5_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_5_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_first = fifof_5_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_first = fifof_5_EMPTY_N ;

  // rule RL_empty_fifof_to_rxe_6_connect_notEmpty
  assign CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_notEmpty = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_notEmpty = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_6_connect_rdy
  assign CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_6_connect_first
  assign CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_first = fifof_6_EMPTY_N ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_first = fifof_6_EMPTY_N ;

  // rule RL_mkConnectionGetPut
  assign CAN_FIRE_RL_mkConnectionGetPut =
	     stage1_RDY_commit_rd_put && stage3_RDY_commit_rd_get ;
  assign WILL_FIRE_RL_mkConnectionGetPut = CAN_FIRE_RL_mkConnectionGetPut ;

  // rule RL_mkConnectionGetPut_1
  assign CAN_FIRE_RL_mkConnectionGetPut_1 = 1'd1 ;
  assign WILL_FIRE_RL_mkConnectionGetPut_1 = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_3_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_ena =
	     fifof_3_EMPTY_N && stage3_rx_stage3_common_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_3_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_ena ;

  // rule RL_empty_txe_to_fifof_3_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_3_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_3_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_3_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_3_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_3_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_4_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_ena =
	     fifof_4_EMPTY_N && stage3_rx_stage3_type_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_4_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_ena ;

  // rule RL_empty_txe_to_fifof_4_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_4_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_4_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_4_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_4_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_4_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_6_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_ena =
	     fifof_6_EMPTY_N && stage3_rx_stage3_dump_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_6_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_ena ;

  // rule RL_empty_txe_to_fifof_6_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_6_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_6_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_6_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_6_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_6_connect_rdy = 1'd1 ;

  // rule RL_gen_new_pc
  assign CAN_FIRE_RL_gen_new_pc =
	     stage3_flush_snd || stage2_mv_redirection_snd ;
  assign WILL_FIRE_RL_gen_new_pc = CAN_FIRE_RL_gen_new_pc ;

  // rule RL_empty_fifof_to_rxe_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_connect_ena =
	     fifof_EMPTY_N && stage2_rx_stage1_operands_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_connect_ena ;

  // rule RL_empty_txe_to_fifof_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_1_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_ena =
	     fifof_1_EMPTY_N && stage2_rx_stage1_control_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_1_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_ena ;

  // rule RL_empty_txe_to_fifof_1_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_1_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_1_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_1_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_1_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_1_connect_rdy = 1'd1 ;

  // rule RL_empty_fifof_to_rxe_2_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_ena =
	     fifof_2_EMPTY_N && stage2_rx_stage1_meta_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_2_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_ena ;

  // rule RL_empty_txe_to_fifof_2_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_2_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_2_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_2_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_2_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_2_connect_rdy = 1'd1 ;

  // rule RL_empty_txe_to_fifof_3_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data =
	     fifof_3_FULL_N && stage2_tx_stage3_common_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data ;

  // rule RL_empty_txe_to_fifof_4_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data =
	     fifof_4_FULL_N && stage2_tx_stage3_type_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data ;

  // rule RL_empty_fifof_to_rxe_5_connect_ena
  assign CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_ena =
	     fifof_5_EMPTY_N && stage2_rx_stage1_dump_deq_ena ;
  assign WILL_FIRE_RL_empty_fifof_to_rxe_5_connect_ena =
	     CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_ena ;

  // rule RL_empty_txe_to_fifof_5_connect_notFull
  assign CAN_FIRE_RL_empty_txe_to_fifof_5_connect_notFull = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_5_connect_notFull = 1'd1 ;

  // rule RL_empty_txe_to_fifof_5_connect_rdy
  assign CAN_FIRE_RL_empty_txe_to_fifof_5_connect_rdy = 1'd1 ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_5_connect_rdy = 1'd1 ;

  // rule RL_redirection_from_stage2
  assign CAN_FIRE_RL_redirection_from_stage2 = stage2_mv_redirection_snd ;
  assign WILL_FIRE_RL_redirection_from_stage2 = stage2_mv_redirection_snd ;

  // rule RL_flush_from_writeback
  assign CAN_FIRE_RL_flush_from_writeback = stage3_flush_snd ;
  assign WILL_FIRE_RL_flush_from_writeback = stage3_flush_snd ;

  // rule RL_empty_txe_to_fifof_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_connect_ena_data =
	     fifof_FULL_N && stage1_tx_stage1_operands_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_connect_ena_data ;

  // rule RL_empty_txe_to_fifof_1_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data =
	     fifof_1_FULL_N && stage1_tx_stage1_control_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data ;

  // rule RL_empty_txe_to_fifof_2_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data =
	     fifof_2_FULL_N && stage1_tx_stage1_meta_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data ;

  // rule RL_empty_txe_to_fifof_5_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data =
	     fifof_5_FULL_N && stage1_tx_stage1_dump_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data ;

  // rule RL_empty_txe_to_fifof_6_connect_ena_data
  assign CAN_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data =
	     fifof_6_FULL_N && stage2_tx_stage3_dump_enq_ena ;
  assign WILL_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data =
	     CAN_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data ;

  // submodule fifof
  assign fifof_D_IN = stage1_tx_stage1_operands_enq_data ;
  assign fifof_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_connect_ena_data ;
  assign fifof_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_connect_ena ;
  assign fifof_CLR = 1'b0 ;

  // submodule fifof_1
  assign fifof_1_D_IN = stage1_tx_stage1_control_enq_data ;
  assign fifof_1_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_1_connect_ena_data ;
  assign fifof_1_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_1_connect_ena ;
  assign fifof_1_CLR = 1'b0 ;

  // submodule fifof_2
  assign fifof_2_D_IN =
	     { stage1_tx_stage1_meta_enq_data[64:43],
	       CASE_stage1tx_stage1_meta_enq_data_BITS_42_TO_ETC__q2,
	       stage1_tx_stage1_meta_enq_data[40:0] } ;
  assign fifof_2_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_2_connect_ena_data ;
  assign fifof_2_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_2_connect_ena ;
  assign fifof_2_CLR = 1'b0 ;

  // submodule fifof_3
  assign fifof_3_D_IN = stage2_tx_stage3_common_enq_data ;
  assign fifof_3_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_3_connect_ena_data ;
  assign fifof_3_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_3_connect_ena ;
  assign fifof_3_CLR = 1'b0 ;

  // submodule fifof_4
  assign fifof_4_D_IN =
	     { CASE_stage2tx_stage3_type_enq_data_BITS_82_TO_ETC__q3,
	       (stage2_tx_stage3_type_enq_data[82:81] == 2'd0) ?
		 { 13'b0101010101010 /* unspecified value */ ,
		   CASE_stage2tx_stage3_type_enq_data_BITS_67_TO_ETC__q4,
		   stage2_tx_stage3_type_enq_data[65:0] } :
		 stage2_tx_stage3_type_enq_data[80:0] } ;
  assign fifof_4_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_4_connect_ena_data ;
  assign fifof_4_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_4_connect_ena ;
  assign fifof_4_CLR = 1'b0 ;

  // submodule fifof_5
  assign fifof_5_D_IN = stage1_tx_stage1_dump_enq_data ;
  assign fifof_5_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_5_connect_ena_data ;
  assign fifof_5_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_5_connect_ena ;
  assign fifof_5_CLR = 1'b0 ;

  // submodule fifof_6
  assign fifof_6_D_IN = stage2_tx_stage3_dump_enq_data ;
  assign fifof_6_ENQ = CAN_FIRE_RL_empty_txe_to_fifof_6_connect_ena_data ;
  assign fifof_6_DEQ = CAN_FIRE_RL_empty_fifof_to_rxe_6_connect_ena ;
  assign fifof_6_CLR = 1'b0 ;

  // submodule stage1
  assign stage1_commit_rd_put = stage3_commit_rd_get ;
  assign stage1_inst_response_put = inst_response_put ;
  assign stage1_ma_csr_decode_c =
	     { (stage3_mv_csr_decode[151:150] == 2'd3) ?
		 stage3_mv_csr_decode[151:150] :
		 2'd0,
	       stage3_mv_csr_decode[149:0] } ;
  assign stage1_ma_csr_misa_c_c = stage3_mv_csr_misa_c ;
  assign stage1_ma_flush_newpc =
	     stage3_flush_snd ? stage3_flush_fst : stage2_mv_redirection_fst ;
  assign stage1_ma_interrupt_i = stage3_mv_interrupt ;
  assign stage1_ma_trigger_data1_t =
	     { CASE_stage3mv_trigger_data1_BITS_43_TO_42_0_s_ETC__q5,
	       CASE_stage3mv_trigger_data1_BITS_21_TO_20_0_s_ETC__q6 } ;
  assign stage1_ma_trigger_data2_t = stage3_mv_trigger_data2 ;
  assign stage1_ma_trigger_enable_t = stage3_mv_trigger_enable ;
  assign stage1_tx_stage1_control_enq_rdy_b = fifof_1_FULL_N ;
  assign stage1_tx_stage1_control_notFull_b = fifof_1_FULL_N ;
  assign stage1_tx_stage1_dump_enq_rdy_b = fifof_5_FULL_N ;
  assign stage1_tx_stage1_dump_notFull_b = fifof_5_FULL_N ;
  assign stage1_tx_stage1_meta_enq_rdy_b = fifof_2_FULL_N ;
  assign stage1_tx_stage1_meta_notFull_b = fifof_2_FULL_N ;
  assign stage1_tx_stage1_operands_enq_rdy_b = fifof_FULL_N ;
  assign stage1_tx_stage1_operands_notFull_b = fifof_FULL_N ;
  assign stage1_EN_inst_request_get = EN_inst_request_get ;
  assign stage1_EN_inst_response_put = EN_inst_response_put ;
  assign stage1_EN_commit_rd_put = CAN_FIRE_RL_mkConnectionGetPut ;
  assign stage1_EN_ma_flush = CAN_FIRE_RL_gen_new_pc ;
  assign stage1_EN_ma_update_eEpoch = stage2_mv_redirection_snd ;
  assign stage1_EN_ma_update_wEpoch = stage3_flush_snd ;

  // submodule stage2
  assign stage2_ma_csr_misa_c_c = stage3_mv_csr_misa_c ;
  assign stage2_ma_trigger_data1_t =
	     { CASE_stage3mv_trigger_data1_BITS_43_TO_42_0_s_ETC__q5,
	       CASE_stage3mv_trigger_data1_BITS_21_TO_20_0_s_ETC__q6 } ;
  assign stage2_ma_trigger_data2_t = stage3_mv_trigger_data2 ;
  assign stage2_ma_trigger_enable_t = stage3_mv_trigger_enable ;
  assign stage2_operand_fwding_put = stage3_operand_fwding_get ;
  assign stage2_rx_stage1_control_first_deq_rdy_b = fifof_1_EMPTY_N ;
  assign stage2_rx_stage1_control_first_x = fifof_1_D_OUT ;
  assign stage2_rx_stage1_control_notEmpty_b = fifof_1_EMPTY_N ;
  assign stage2_rx_stage1_dump_first_deq_rdy_b = fifof_5_EMPTY_N ;
  assign stage2_rx_stage1_dump_first_x = fifof_5_D_OUT ;
  assign stage2_rx_stage1_dump_notEmpty_b = fifof_5_EMPTY_N ;
  assign stage2_rx_stage1_meta_first_deq_rdy_b = fifof_2_EMPTY_N ;
  assign stage2_rx_stage1_meta_first_x =
	     { fifof_2_D_OUT[64:43],
	       CASE_IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_fi_ETC__q7,
	       fifof_2_D_OUT[40:0] } ;
  assign stage2_rx_stage1_meta_notEmpty_b = fifof_2_EMPTY_N ;
  assign stage2_rx_stage1_operands_first_deq_rdy_b = fifof_EMPTY_N ;
  assign stage2_rx_stage1_operands_first_x = fifof_D_OUT ;
  assign stage2_rx_stage1_operands_notEmpty_b = fifof_EMPTY_N ;
  assign stage2_tx_stage3_common_enq_rdy_b = fifof_3_FULL_N ;
  assign stage2_tx_stage3_common_notFull_b = fifof_3_FULL_N ;
  assign stage2_tx_stage3_dump_enq_rdy_b = fifof_6_FULL_N ;
  assign stage2_tx_stage3_dump_notFull_b = fifof_6_FULL_N ;
  assign stage2_tx_stage3_type_enq_rdy_b = fifof_4_FULL_N ;
  assign stage2_tx_stage3_type_notFull_b = fifof_4_FULL_N ;
  assign stage2_EN_memory_request_get = EN_memory_request_get ;
  assign stage2_EN_operand_fwding_put = 1'd1 ;
  assign stage2_EN_ma_update_wEpoch = stage3_flush_snd ;
  assign stage2_EN_ma_csr_misa_c = 1'd1 ;

  // submodule stage3
  assign stage3_clint_msip_intrpt = clint_msip_intrpt ;
  assign stage3_clint_mtime_c_mtime = clint_mtime_c_mtime ;
  assign stage3_clint_mtip_intrpt = clint_mtip_intrpt ;
  assign stage3_ext_interrupt_i = ext_interrupt_intrpt ;
  assign stage3_ma_delayed_output_r = stage2_mv_delayed_output ;
  assign stage3_memory_response_put = memory_response_put ;
  assign stage3_rx_stage3_common_first_deq_rdy_b = fifof_3_EMPTY_N ;
  assign stage3_rx_stage3_common_first_x = fifof_3_D_OUT ;
  assign stage3_rx_stage3_common_notEmpty_b = fifof_3_EMPTY_N ;
  assign stage3_rx_stage3_dump_first_deq_rdy_b = fifof_6_EMPTY_N ;
  assign stage3_rx_stage3_dump_first_x = fifof_6_D_OUT ;
  assign stage3_rx_stage3_dump_notEmpty_b = fifof_6_EMPTY_N ;
  assign stage3_rx_stage3_type_first_deq_rdy_b = fifof_4_EMPTY_N ;
  assign stage3_rx_stage3_type_first_x =
	     (fifof_4_EMPTY_N && fifof_4_D_OUT[82:81] == 2'd0) ?
	       { 2'd0,
		 13'b0101010101010 /* unspecified value */ ,
		 CASE_IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_f_ETC__q8,
		 fifof_4_D_OUT[65:0] } :
	       { (fifof_4_EMPTY_N && fifof_4_D_OUT[82:81] == 2'd1) ?
		   2'd1 :
		   ((fifof_4_EMPTY_N && fifof_4_D_OUT[82:81] == 2'd2) ?
		      2'd2 :
		      2'd3),
		 fifof_4_D_OUT[80:0] } ;
  assign stage3_rx_stage3_type_notEmpty_b = fifof_4_EMPTY_N ;
  assign stage3_EN_memory_response_put = EN_memory_response_put ;
  assign stage3_EN_commit_rd_get = CAN_FIRE_RL_mkConnectionGetPut ;
  assign stage3_EN_operand_fwding_get = 1'd1 ;
  assign stage3_EN_clint_msip = EN_clint_msip ;
  assign stage3_EN_clint_mtip = EN_clint_mtip ;
  assign stage3_EN_clint_mtime = EN_clint_mtime ;
  assign stage3_EN_ext_interrupt = EN_ext_interrupt ;
  assign stage3_EN_dump_get = EN_dump_get ;
  assign stage3_EN_ma_delayed_output = 1'd1 ;

  // remaining internal signals
  always@(stage2_memory_request_get)
  begin
    case (stage2_memory_request_get[10:9])
      2'd0, 2'd1, 2'd3:
	  CASE_stage2memory_request_get_BITS_10_TO_9_0__ETC__q1 =
	      stage2_memory_request_get[10:9];
      2'd2: CASE_stage2memory_request_get_BITS_10_TO_9_0__ETC__q1 = 2'd2;
    endcase
  end
  always@(fifof_2_D_OUT)
  begin
    case (fifof_2_D_OUT[42:41])
      2'd0, 2'd1:
	  IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57 =
	      fifof_2_D_OUT[42:41];
      2'd2: IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57 = 2'd3;
      2'd3: IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57 = 2'd2;
    endcase
  end
  always@(fifof_4_D_OUT)
  begin
    case (fifof_4_D_OUT[67:66])
      2'd0, 2'd1:
	  IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121 =
	      fifof_4_D_OUT[67:66];
      2'd2: IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121 = 2'd3;
      2'd3: IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121 = 2'd2;
    endcase
  end
  always@(stage1_tx_stage1_meta_enq_data)
  begin
    case (stage1_tx_stage1_meta_enq_data[42:41])
      2'd0, 2'd1, 2'd3:
	  CASE_stage1tx_stage1_meta_enq_data_BITS_42_TO_ETC__q2 =
	      stage1_tx_stage1_meta_enq_data[42:41];
      2'd2: CASE_stage1tx_stage1_meta_enq_data_BITS_42_TO_ETC__q2 = 2'd2;
    endcase
  end
  always@(stage2_tx_stage3_type_enq_data)
  begin
    case (stage2_tx_stage3_type_enq_data[82:81])
      2'd0, 2'd1, 2'd2:
	  CASE_stage2tx_stage3_type_enq_data_BITS_82_TO_ETC__q3 =
	      stage2_tx_stage3_type_enq_data[82:81];
      2'd3: CASE_stage2tx_stage3_type_enq_data_BITS_82_TO_ETC__q3 = 2'd3;
    endcase
  end
  always@(stage2_tx_stage3_type_enq_data)
  begin
    case (stage2_tx_stage3_type_enq_data[67:66])
      2'd0, 2'd1, 2'd3:
	  CASE_stage2tx_stage3_type_enq_data_BITS_67_TO_ETC__q4 =
	      stage2_tx_stage3_type_enq_data[67:66];
      2'd2: CASE_stage2tx_stage3_type_enq_data_BITS_67_TO_ETC__q4 = 2'd2;
    endcase
  end
  always@(stage3_mv_trigger_data1)
  begin
    case (stage3_mv_trigger_data1[43:42])
      2'd0, 2'd1, 2'd2:
	  CASE_stage3mv_trigger_data1_BITS_43_TO_42_0_s_ETC__q5 =
	      stage3_mv_trigger_data1[43:22];
      2'd3:
	  CASE_stage3mv_trigger_data1_BITS_43_TO_42_0_s_ETC__q5 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(stage3_mv_trigger_data1)
  begin
    case (stage3_mv_trigger_data1[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_stage3mv_trigger_data1_BITS_21_TO_20_0_s_ETC__q6 =
	      stage3_mv_trigger_data1[21:0];
      2'd3:
	  CASE_stage3mv_trigger_data1_BITS_21_TO_20_0_s_ETC__q6 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57)
  begin
    case (IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57)
      2'd0, 2'd1:
	  CASE_IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_fi_ETC__q7 =
	      IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_first___ETC___d57;
      2'd2: CASE_IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_fi_ETC__q7 = 2'd3;
      2'd3: CASE_IF_fifof_2_notEmpty__1_THEN_IF_fifof_2_fi_ETC__q7 = 2'd2;
    endcase
  end
  always@(IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121)
  begin
    case (IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121)
      2'd0, 2'd1:
	  CASE_IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_f_ETC__q8 =
	      IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_first__ETC___d121;
      2'd2: CASE_IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_f_ETC__q8 = 2'd3;
      2'd3: CASE_IF_fifof_4_notEmpty__08_THEN_IF_fifof_4_f_ETC__q8 = 2'd2;
    endcase
  end
endmodule  // mkriscv

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:52 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// master_awvalid                 O     1 reg
// master_awaddr                  O    32 reg
// master_awprot                  O     3 reg
// master_awsize                  O     2 reg
// master_wvalid                  O     1 reg
// master_wdata                   O    64 reg
// master_wstrb                   O     8 reg
// master_bready                  O     1 reg
// master_arvalid                 O     1 reg
// master_araddr                  O    32 reg
// master_arprot                  O     3 reg
// master_arsize                  O     2 reg
// master_rready                  O     1 reg
// slave_awready                  O     1 reg
// slave_wready                   O     1 reg
// slave_bvalid                   O     1 reg
// slave_bresp                    O     2 reg
// slave_arready                  O     1 reg
// slave_rvalid                   O     1 reg
// slave_rresp                    O     2 reg
// slave_rdata                    O    64 reg
// mv_end_simulation              O     1
// RDY_mv_end_simulation          O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// master_m_awready_awready       I     1
// master_m_wready_wready         I     1
// master_m_bvalid_bvalid         I     1
// master_m_bvalid_bresp          I     2 reg
// master_m_arready_arready       I     1
// master_m_rvalid_rvalid         I     1
// master_m_rvalid_rresp          I     2 reg
// master_m_rvalid_rdata          I    64 reg
// slave_m_awvalid_awvalid        I     1
// slave_m_awvalid_awaddr         I    32 reg
// slave_m_awvalid_awsize         I     2 reg
// slave_m_awvalid_awprot         I     3 reg
// slave_m_wvalid_wvalid          I     1
// slave_m_wvalid_wdata           I    64 reg
// slave_m_wvalid_wstrb           I     8 reg
// slave_m_bready_bready          I     1
// slave_m_arvalid_arvalid        I     1
// slave_m_arvalid_araddr         I    32 reg
// slave_m_arvalid_arsize         I     2 reg
// slave_m_arvalid_arprot         I     3 reg
// slave_m_rready_rready          I     1
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mksign_dump_axi4lite(CLK,
			    RST_N,

			    master_awvalid,

			    master_awaddr,

			    master_awprot,

			    master_awsize,

			    master_m_awready_awready,

			    master_wvalid,

			    master_wdata,

			    master_wstrb,

			    master_m_wready_wready,

			    master_m_bvalid_bvalid,
			    master_m_bvalid_bresp,

			    master_bready,

			    master_arvalid,

			    master_araddr,

			    master_arprot,

			    master_arsize,

			    master_m_arready_arready,

			    master_m_rvalid_rvalid,
			    master_m_rvalid_rresp,
			    master_m_rvalid_rdata,

			    master_rready,

			    slave_m_awvalid_awvalid,
			    slave_m_awvalid_awaddr,
			    slave_m_awvalid_awsize,
			    slave_m_awvalid_awprot,

			    slave_awready,

			    slave_m_wvalid_wvalid,
			    slave_m_wvalid_wdata,
			    slave_m_wvalid_wstrb,

			    slave_wready,

			    slave_bvalid,

			    slave_bresp,

			    slave_m_bready_bready,

			    slave_m_arvalid_arvalid,
			    slave_m_arvalid_araddr,
			    slave_m_arvalid_arsize,
			    slave_m_arvalid_arprot,

			    slave_arready,

			    slave_rvalid,

			    slave_rresp,

			    slave_rdata,

			    slave_m_rready_rready,

			    mv_end_simulation,
			    RDY_mv_end_simulation);
  input  CLK;
  input  RST_N;

  // value method master_m_awvalid
  output master_awvalid;

  // value method master_m_awaddr
  output [31 : 0] master_awaddr;

  // value method master_m_awuser

  // value method master_m_awprot
  output [2 : 0] master_awprot;

  // value method master_m_awsize
  output [1 : 0] master_awsize;

  // action method master_m_awready
  input  master_m_awready_awready;

  // value method master_m_wvalid
  output master_wvalid;

  // value method master_m_wdata
  output [63 : 0] master_wdata;

  // value method master_m_wstrb
  output [7 : 0] master_wstrb;

  // action method master_m_wready
  input  master_m_wready_wready;

  // action method master_m_bvalid
  input  master_m_bvalid_bvalid;
  input  [1 : 0] master_m_bvalid_bresp;

  // value method master_m_bready
  output master_bready;

  // value method master_m_arvalid
  output master_arvalid;

  // value method master_m_araddr
  output [31 : 0] master_araddr;

  // value method master_m_aruser

  // value method master_m_arprot
  output [2 : 0] master_arprot;

  // value method master_m_arsize
  output [1 : 0] master_arsize;

  // action method master_m_arready
  input  master_m_arready_arready;

  // action method master_m_rvalid
  input  master_m_rvalid_rvalid;
  input  [1 : 0] master_m_rvalid_rresp;
  input  [63 : 0] master_m_rvalid_rdata;

  // value method master_m_rready
  output master_rready;

  // action method slave_m_awvalid
  input  slave_m_awvalid_awvalid;
  input  [31 : 0] slave_m_awvalid_awaddr;
  input  [1 : 0] slave_m_awvalid_awsize;
  input  [2 : 0] slave_m_awvalid_awprot;

  // value method slave_m_awready
  output slave_awready;

  // action method slave_m_wvalid
  input  slave_m_wvalid_wvalid;
  input  [63 : 0] slave_m_wvalid_wdata;
  input  [7 : 0] slave_m_wvalid_wstrb;

  // value method slave_m_wready
  output slave_wready;

  // value method slave_m_bvalid
  output slave_bvalid;

  // value method slave_m_bresp
  output [1 : 0] slave_bresp;

  // value method slave_m_buser

  // action method slave_m_bready
  input  slave_m_bready_bready;

  // action method slave_m_arvalid
  input  slave_m_arvalid_arvalid;
  input  [31 : 0] slave_m_arvalid_araddr;
  input  [1 : 0] slave_m_arvalid_arsize;
  input  [2 : 0] slave_m_arvalid_arprot;

  // value method slave_m_arready
  output slave_arready;

  // value method slave_m_rvalid
  output slave_rvalid;

  // value method slave_m_rresp
  output [1 : 0] slave_rresp;

  // value method slave_m_rdata
  output [63 : 0] slave_rdata;

  // value method slave_m_ruser

  // action method slave_m_rready
  input  slave_m_rready_rready;

  // value method mv_end_simulation
  output mv_end_simulation;
  output RDY_mv_end_simulation;

  // signals for module outputs
  wire [63 : 0] master_wdata, slave_rdata;
  wire [31 : 0] master_araddr, master_awaddr;
  wire [7 : 0] master_wstrb;
  wire [2 : 0] master_arprot, master_awprot;
  wire [1 : 0] master_arsize, master_awsize, slave_bresp, slave_rresp;
  wire RDY_mv_end_simulation,
       master_arvalid,
       master_awvalid,
       master_bready,
       master_rready,
       master_wvalid,
       mv_end_simulation,
       slave_arready,
       slave_awready,
       slave_bvalid,
       slave_rvalid,
       slave_wready;

  // inlined wires
  wire rg_end_sim_EN_port0__write, rg_end_sim_port1__read;

  // register dataarray_0
  reg [31 : 0] dataarray_0;
  wire [31 : 0] dataarray_0_D_IN;
  wire dataarray_0_EN;

  // register dataarray_1
  reg [31 : 0] dataarray_1;
  wire [31 : 0] dataarray_1_D_IN;
  wire dataarray_1_EN;

  // register dump
  reg [31 : 0] dump;
  wire [31 : 0] dump_D_IN;
  wire dump_EN;

  // register rg_cnt
  reg [4 : 0] rg_cnt;
  wire [4 : 0] rg_cnt_D_IN;
  wire rg_cnt_EN;

  // register rg_end_address
  reg [31 : 0] rg_end_address;
  wire [31 : 0] rg_end_address_D_IN;
  wire rg_end_address_EN;

  // register rg_end_sim
  reg rg_end_sim;
  wire rg_end_sim_D_IN, rg_end_sim_EN;

  // register rg_start
  reg rg_start;
  wire rg_start_D_IN, rg_start_EN;

  // register rg_start_address
  reg [31 : 0] rg_start_address;
  wire [31 : 0] rg_start_address_D_IN;
  wire rg_start_address_EN;

  // register rg_total_count
  reg [31 : 0] rg_total_count;
  wire [31 : 0] rg_total_count_D_IN;
  wire rg_total_count_EN;

  // register rg_word_count
  reg rg_word_count;
  wire rg_word_count_D_IN, rg_word_count_EN;

  // ports of submodule ff_lower_order_bits
  wire [2 : 0] ff_lower_order_bits_D_IN, ff_lower_order_bits_D_OUT;
  wire ff_lower_order_bits_CLR,
       ff_lower_order_bits_DEQ,
       ff_lower_order_bits_EMPTY_N,
       ff_lower_order_bits_ENQ,
       ff_lower_order_bits_FULL_N;

  // ports of submodule m_xactor_f_rd_addr
  wire [36 : 0] m_xactor_f_rd_addr_D_IN, m_xactor_f_rd_addr_D_OUT;
  wire m_xactor_f_rd_addr_CLR,
       m_xactor_f_rd_addr_DEQ,
       m_xactor_f_rd_addr_EMPTY_N,
       m_xactor_f_rd_addr_ENQ,
       m_xactor_f_rd_addr_FULL_N;

  // ports of submodule m_xactor_f_rd_data
  wire [65 : 0] m_xactor_f_rd_data_D_IN, m_xactor_f_rd_data_D_OUT;
  wire m_xactor_f_rd_data_CLR,
       m_xactor_f_rd_data_DEQ,
       m_xactor_f_rd_data_EMPTY_N,
       m_xactor_f_rd_data_ENQ,
       m_xactor_f_rd_data_FULL_N;

  // ports of submodule m_xactor_f_wr_addr
  wire [36 : 0] m_xactor_f_wr_addr_D_IN, m_xactor_f_wr_addr_D_OUT;
  wire m_xactor_f_wr_addr_CLR,
       m_xactor_f_wr_addr_DEQ,
       m_xactor_f_wr_addr_EMPTY_N,
       m_xactor_f_wr_addr_ENQ;

  // ports of submodule m_xactor_f_wr_data
  wire [71 : 0] m_xactor_f_wr_data_D_IN, m_xactor_f_wr_data_D_OUT;
  wire m_xactor_f_wr_data_CLR,
       m_xactor_f_wr_data_DEQ,
       m_xactor_f_wr_data_EMPTY_N,
       m_xactor_f_wr_data_ENQ;

  // ports of submodule m_xactor_f_wr_resp
  wire [1 : 0] m_xactor_f_wr_resp_D_IN;
  wire m_xactor_f_wr_resp_CLR,
       m_xactor_f_wr_resp_DEQ,
       m_xactor_f_wr_resp_ENQ,
       m_xactor_f_wr_resp_FULL_N;

  // ports of submodule s_xactor_f_rd_addr
  wire [36 : 0] s_xactor_f_rd_addr_D_IN;
  wire s_xactor_f_rd_addr_CLR,
       s_xactor_f_rd_addr_DEQ,
       s_xactor_f_rd_addr_ENQ,
       s_xactor_f_rd_addr_FULL_N;

  // ports of submodule s_xactor_f_rd_data
  wire [65 : 0] s_xactor_f_rd_data_D_IN, s_xactor_f_rd_data_D_OUT;
  wire s_xactor_f_rd_data_CLR,
       s_xactor_f_rd_data_DEQ,
       s_xactor_f_rd_data_EMPTY_N,
       s_xactor_f_rd_data_ENQ;

  // ports of submodule s_xactor_f_wr_addr
  wire [36 : 0] s_xactor_f_wr_addr_D_IN, s_xactor_f_wr_addr_D_OUT;
  wire s_xactor_f_wr_addr_CLR,
       s_xactor_f_wr_addr_DEQ,
       s_xactor_f_wr_addr_EMPTY_N,
       s_xactor_f_wr_addr_ENQ,
       s_xactor_f_wr_addr_FULL_N;

  // ports of submodule s_xactor_f_wr_data
  wire [71 : 0] s_xactor_f_wr_data_D_IN, s_xactor_f_wr_data_D_OUT;
  wire s_xactor_f_wr_data_CLR,
       s_xactor_f_wr_data_DEQ,
       s_xactor_f_wr_data_EMPTY_N,
       s_xactor_f_wr_data_ENQ,
       s_xactor_f_wr_data_FULL_N;

  // ports of submodule s_xactor_f_wr_resp
  reg [1 : 0] s_xactor_f_wr_resp_D_IN;
  wire [1 : 0] s_xactor_f_wr_resp_D_OUT;
  wire s_xactor_f_wr_resp_CLR,
       s_xactor_f_wr_resp_DEQ,
       s_xactor_f_wr_resp_EMPTY_N,
       s_xactor_f_wr_resp_ENQ,
       s_xactor_f_wr_resp_FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_configure_registers,
       CAN_FIRE_RL_open_file,
       CAN_FIRE_RL_receive_response,
       CAN_FIRE_RL_send_request,
       CAN_FIRE_master_m_arready,
       CAN_FIRE_master_m_awready,
       CAN_FIRE_master_m_bvalid,
       CAN_FIRE_master_m_rvalid,
       CAN_FIRE_master_m_wready,
       CAN_FIRE_slave_m_arvalid,
       CAN_FIRE_slave_m_awvalid,
       CAN_FIRE_slave_m_bready,
       CAN_FIRE_slave_m_rready,
       CAN_FIRE_slave_m_wvalid,
       WILL_FIRE_RL_configure_registers,
       WILL_FIRE_RL_open_file,
       WILL_FIRE_RL_receive_response,
       WILL_FIRE_RL_send_request,
       WILL_FIRE_master_m_arready,
       WILL_FIRE_master_m_awready,
       WILL_FIRE_master_m_bvalid,
       WILL_FIRE_master_m_rvalid,
       WILL_FIRE_master_m_wready,
       WILL_FIRE_slave_m_arvalid,
       WILL_FIRE_slave_m_awvalid,
       WILL_FIRE_slave_m_bready,
       WILL_FIRE_slave_m_rready,
       WILL_FIRE_slave_m_wvalid;

  // inputs to muxes for submodule ports
  wire [31 : 0] MUX_rg_start_address_write_1__VAL_2,
		MUX_rg_total_count_write_1__VAL_1,
		MUX_rg_total_count_write_1__VAL_2;
  wire MUX_rg_start_write_1__SEL_1,
       MUX_rg_start_address_write_1__SEL_1,
       MUX_rg_start_address_write_1__SEL_2,
       MUX_rg_total_count_write_1__SEL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg [31 : 0] TASK_fopen___d3;
  reg [63 : 0] v__h2897;
  // synopsys translate_on

  // remaining internal signals
  wire [63 : 0] m_xactor_f_rd_dataD_OUT_BITS_63_TO_0_SRL_lv_s_ETC__q2;
  wire [31 : 0] s_xactor_f_wr_dataD_OUT_BITS_39_TO_8_MINUS_rg_ETC__q1;
  wire [5 : 0] lv_shift__h2655;
  wire rg_cnt_ULT_5___d2, rg_start_address_0_ULT_rg_end_address_4___d35;

  // value method master_m_awvalid
  assign master_awvalid = m_xactor_f_wr_addr_EMPTY_N ;

  // value method master_m_awaddr
  assign master_awaddr = m_xactor_f_wr_addr_D_OUT[36:5] ;

  // value method master_m_awprot
  assign master_awprot = m_xactor_f_wr_addr_D_OUT[4:2] ;

  // value method master_m_awsize
  assign master_awsize = m_xactor_f_wr_addr_D_OUT[1:0] ;

  // action method master_m_awready
  assign CAN_FIRE_master_m_awready = 1'd1 ;
  assign WILL_FIRE_master_m_awready = 1'd1 ;

  // value method master_m_wvalid
  assign master_wvalid = m_xactor_f_wr_data_EMPTY_N ;

  // value method master_m_wdata
  assign master_wdata = m_xactor_f_wr_data_D_OUT[71:8] ;

  // value method master_m_wstrb
  assign master_wstrb = m_xactor_f_wr_data_D_OUT[7:0] ;

  // action method master_m_wready
  assign CAN_FIRE_master_m_wready = 1'd1 ;
  assign WILL_FIRE_master_m_wready = 1'd1 ;

  // action method master_m_bvalid
  assign CAN_FIRE_master_m_bvalid = 1'd1 ;
  assign WILL_FIRE_master_m_bvalid = 1'd1 ;

  // value method master_m_bready
  assign master_bready = m_xactor_f_wr_resp_FULL_N ;

  // value method master_m_arvalid
  assign master_arvalid = m_xactor_f_rd_addr_EMPTY_N ;

  // value method master_m_araddr
  assign master_araddr = m_xactor_f_rd_addr_D_OUT[36:5] ;

  // value method master_m_arprot
  assign master_arprot = m_xactor_f_rd_addr_D_OUT[4:2] ;

  // value method master_m_arsize
  assign master_arsize = m_xactor_f_rd_addr_D_OUT[1:0] ;

  // action method master_m_arready
  assign CAN_FIRE_master_m_arready = 1'd1 ;
  assign WILL_FIRE_master_m_arready = 1'd1 ;

  // action method master_m_rvalid
  assign CAN_FIRE_master_m_rvalid = 1'd1 ;
  assign WILL_FIRE_master_m_rvalid = 1'd1 ;

  // value method master_m_rready
  assign master_rready = m_xactor_f_rd_data_FULL_N ;

  // action method slave_m_awvalid
  assign CAN_FIRE_slave_m_awvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_awvalid = 1'd1 ;

  // value method slave_m_awready
  assign slave_awready = s_xactor_f_wr_addr_FULL_N ;

  // action method slave_m_wvalid
  assign CAN_FIRE_slave_m_wvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_wvalid = 1'd1 ;

  // value method slave_m_wready
  assign slave_wready = s_xactor_f_wr_data_FULL_N ;

  // value method slave_m_bvalid
  assign slave_bvalid = s_xactor_f_wr_resp_EMPTY_N ;

  // value method slave_m_bresp
  assign slave_bresp = s_xactor_f_wr_resp_D_OUT ;

  // action method slave_m_bready
  assign CAN_FIRE_slave_m_bready = 1'd1 ;
  assign WILL_FIRE_slave_m_bready = 1'd1 ;

  // action method slave_m_arvalid
  assign CAN_FIRE_slave_m_arvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_arvalid = 1'd1 ;

  // value method slave_m_arready
  assign slave_arready = s_xactor_f_rd_addr_FULL_N ;

  // value method slave_m_rvalid
  assign slave_rvalid = s_xactor_f_rd_data_EMPTY_N ;

  // value method slave_m_rresp
  assign slave_rresp = s_xactor_f_rd_data_D_OUT[65:64] ;

  // value method slave_m_rdata
  assign slave_rdata = s_xactor_f_rd_data_D_OUT[63:0] ;

  // action method slave_m_rready
  assign CAN_FIRE_slave_m_rready = 1'd1 ;
  assign WILL_FIRE_slave_m_rready = 1'd1 ;

  // value method mv_end_simulation
  assign mv_end_simulation = rg_end_sim_EN_port0__write || rg_end_sim ;
  assign RDY_mv_end_simulation = 1'd1 ;

  // submodule ff_lower_order_bits
  SizedFIFO #(.p1width(32'd3),
	      .p2depth(32'd8),
	      .p3cntr_width(32'd3),
	      .guarded(32'd1)) ff_lower_order_bits(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(ff_lower_order_bits_D_IN),
						   .ENQ(ff_lower_order_bits_ENQ),
						   .DEQ(ff_lower_order_bits_DEQ),
						   .CLR(ff_lower_order_bits_CLR),
						   .D_OUT(ff_lower_order_bits_D_OUT),
						   .FULL_N(ff_lower_order_bits_FULL_N),
						   .EMPTY_N(ff_lower_order_bits_EMPTY_N));

  // submodule m_xactor_f_rd_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) m_xactor_f_rd_addr(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(m_xactor_f_rd_addr_D_IN),
							      .ENQ(m_xactor_f_rd_addr_ENQ),
							      .DEQ(m_xactor_f_rd_addr_DEQ),
							      .CLR(m_xactor_f_rd_addr_CLR),
							      .D_OUT(m_xactor_f_rd_addr_D_OUT),
							      .FULL_N(m_xactor_f_rd_addr_FULL_N),
							      .EMPTY_N(m_xactor_f_rd_addr_EMPTY_N));

  // submodule m_xactor_f_rd_data
  FIFO2 #(.width(32'd66), .guarded(32'd1)) m_xactor_f_rd_data(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(m_xactor_f_rd_data_D_IN),
							      .ENQ(m_xactor_f_rd_data_ENQ),
							      .DEQ(m_xactor_f_rd_data_DEQ),
							      .CLR(m_xactor_f_rd_data_CLR),
							      .D_OUT(m_xactor_f_rd_data_D_OUT),
							      .FULL_N(m_xactor_f_rd_data_FULL_N),
							      .EMPTY_N(m_xactor_f_rd_data_EMPTY_N));

  // submodule m_xactor_f_wr_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) m_xactor_f_wr_addr(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(m_xactor_f_wr_addr_D_IN),
							      .ENQ(m_xactor_f_wr_addr_ENQ),
							      .DEQ(m_xactor_f_wr_addr_DEQ),
							      .CLR(m_xactor_f_wr_addr_CLR),
							      .D_OUT(m_xactor_f_wr_addr_D_OUT),
							      .FULL_N(),
							      .EMPTY_N(m_xactor_f_wr_addr_EMPTY_N));

  // submodule m_xactor_f_wr_data
  FIFO2 #(.width(32'd72), .guarded(32'd1)) m_xactor_f_wr_data(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(m_xactor_f_wr_data_D_IN),
							      .ENQ(m_xactor_f_wr_data_ENQ),
							      .DEQ(m_xactor_f_wr_data_DEQ),
							      .CLR(m_xactor_f_wr_data_CLR),
							      .D_OUT(m_xactor_f_wr_data_D_OUT),
							      .FULL_N(),
							      .EMPTY_N(m_xactor_f_wr_data_EMPTY_N));

  // submodule m_xactor_f_wr_resp
  FIFO2 #(.width(32'd2), .guarded(32'd1)) m_xactor_f_wr_resp(.RST(RST_N),
							     .CLK(CLK),
							     .D_IN(m_xactor_f_wr_resp_D_IN),
							     .ENQ(m_xactor_f_wr_resp_ENQ),
							     .DEQ(m_xactor_f_wr_resp_DEQ),
							     .CLR(m_xactor_f_wr_resp_CLR),
							     .D_OUT(),
							     .FULL_N(m_xactor_f_wr_resp_FULL_N),
							     .EMPTY_N());

  // submodule s_xactor_f_rd_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) s_xactor_f_rd_addr(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(s_xactor_f_rd_addr_D_IN),
							      .ENQ(s_xactor_f_rd_addr_ENQ),
							      .DEQ(s_xactor_f_rd_addr_DEQ),
							      .CLR(s_xactor_f_rd_addr_CLR),
							      .D_OUT(),
							      .FULL_N(s_xactor_f_rd_addr_FULL_N),
							      .EMPTY_N());

  // submodule s_xactor_f_rd_data
  FIFO2 #(.width(32'd66), .guarded(32'd1)) s_xactor_f_rd_data(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(s_xactor_f_rd_data_D_IN),
							      .ENQ(s_xactor_f_rd_data_ENQ),
							      .DEQ(s_xactor_f_rd_data_DEQ),
							      .CLR(s_xactor_f_rd_data_CLR),
							      .D_OUT(s_xactor_f_rd_data_D_OUT),
							      .FULL_N(),
							      .EMPTY_N(s_xactor_f_rd_data_EMPTY_N));

  // submodule s_xactor_f_wr_addr
  FIFO2 #(.width(32'd37), .guarded(32'd1)) s_xactor_f_wr_addr(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(s_xactor_f_wr_addr_D_IN),
							      .ENQ(s_xactor_f_wr_addr_ENQ),
							      .DEQ(s_xactor_f_wr_addr_DEQ),
							      .CLR(s_xactor_f_wr_addr_CLR),
							      .D_OUT(s_xactor_f_wr_addr_D_OUT),
							      .FULL_N(s_xactor_f_wr_addr_FULL_N),
							      .EMPTY_N(s_xactor_f_wr_addr_EMPTY_N));

  // submodule s_xactor_f_wr_data
  FIFO2 #(.width(32'd72), .guarded(32'd1)) s_xactor_f_wr_data(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(s_xactor_f_wr_data_D_IN),
							      .ENQ(s_xactor_f_wr_data_ENQ),
							      .DEQ(s_xactor_f_wr_data_DEQ),
							      .CLR(s_xactor_f_wr_data_CLR),
							      .D_OUT(s_xactor_f_wr_data_D_OUT),
							      .FULL_N(s_xactor_f_wr_data_FULL_N),
							      .EMPTY_N(s_xactor_f_wr_data_EMPTY_N));

  // submodule s_xactor_f_wr_resp
  FIFO2 #(.width(32'd2), .guarded(32'd1)) s_xactor_f_wr_resp(.RST(RST_N),
							     .CLK(CLK),
							     .D_IN(s_xactor_f_wr_resp_D_IN),
							     .ENQ(s_xactor_f_wr_resp_ENQ),
							     .DEQ(s_xactor_f_wr_resp_DEQ),
							     .CLR(s_xactor_f_wr_resp_CLR),
							     .D_OUT(s_xactor_f_wr_resp_D_OUT),
							     .FULL_N(s_xactor_f_wr_resp_FULL_N),
							     .EMPTY_N(s_xactor_f_wr_resp_EMPTY_N));

  // rule RL_open_file
  assign CAN_FIRE_RL_open_file = rg_cnt_ULT_5___d2 ;
  assign WILL_FIRE_RL_open_file = rg_cnt_ULT_5___d2 ;

  // rule RL_configure_registers
  assign CAN_FIRE_RL_configure_registers =
	     s_xactor_f_wr_addr_EMPTY_N && s_xactor_f_wr_data_EMPTY_N &&
	     s_xactor_f_wr_resp_FULL_N &&
	     !rg_start ;
  assign WILL_FIRE_RL_configure_registers = CAN_FIRE_RL_configure_registers ;

  // rule RL_send_request
  assign CAN_FIRE_RL_send_request =
	     m_xactor_f_rd_addr_FULL_N && ff_lower_order_bits_FULL_N &&
	     rg_start ;
  assign WILL_FIRE_RL_send_request = CAN_FIRE_RL_send_request ;

  // rule RL_receive_response
  assign CAN_FIRE_RL_receive_response =
	     m_xactor_f_rd_data_EMPTY_N && ff_lower_order_bits_EMPTY_N &&
	     !rg_cnt_ULT_5___d2 &&
	     rg_start ;
  assign WILL_FIRE_RL_receive_response = CAN_FIRE_RL_receive_response ;

  // inputs to muxes for submodule ports
  assign MUX_rg_start_write_1__SEL_1 =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h8 &&
	     rg_start_address != s_xactor_f_wr_data_D_OUT[39:8] ;
  assign MUX_rg_start_address_write_1__SEL_1 =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h0 ;
  assign MUX_rg_start_address_write_1__SEL_2 =
	     WILL_FIRE_RL_send_request &&
	     rg_start_address_0_ULT_rg_end_address_4___d35 ;
  assign MUX_rg_total_count_write_1__SEL_1 =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h8 ;
  assign MUX_rg_start_address_write_1__VAL_2 = rg_start_address + 32'd4 ;
  assign MUX_rg_total_count_write_1__VAL_1 =
	     { 2'd0,
	       s_xactor_f_wr_dataD_OUT_BITS_39_TO_8_MINUS_rg_ETC__q1[31:2] } ;
  assign MUX_rg_total_count_write_1__VAL_2 = rg_total_count - 32'd1 ;

  // inlined wires
  assign rg_end_sim_EN_port0__write =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'hC ;
  assign rg_end_sim_port1__read = rg_end_sim_EN_port0__write || rg_end_sim ;

  // register dataarray_0
  assign dataarray_0_D_IN = 32'h0 ;
  assign dataarray_0_EN = 1'b0 ;

  // register dataarray_1
  assign dataarray_1_D_IN = 32'h0 ;
  assign dataarray_1_EN = 1'b0 ;

  // register dump
  assign dump_D_IN = TASK_fopen___d3 ;
  assign dump_EN = rg_cnt_ULT_5___d2 ;

  // register rg_cnt
  assign rg_cnt_D_IN = rg_cnt + 5'd1 ;
  assign rg_cnt_EN = rg_cnt_ULT_5___d2 ;

  // register rg_end_address
  assign rg_end_address_D_IN = s_xactor_f_wr_data_D_OUT[39:8] ;
  assign rg_end_address_EN = MUX_rg_total_count_write_1__SEL_1 ;

  // register rg_end_sim
  assign rg_end_sim_D_IN = rg_end_sim_port1__read ;
  assign rg_end_sim_EN = 1'b1 ;

  // register rg_start
  assign rg_start_D_IN = MUX_rg_start_write_1__SEL_1 ;
  assign rg_start_EN =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h8 &&
	     rg_start_address != s_xactor_f_wr_data_D_OUT[39:8] ||
	     WILL_FIRE_RL_receive_response && rg_total_count == 32'd1 ;

  // register rg_start_address
  assign rg_start_address_D_IN =
	     MUX_rg_start_address_write_1__SEL_1 ?
	       s_xactor_f_wr_data_D_OUT[39:8] :
	       MUX_rg_start_address_write_1__VAL_2 ;
  assign rg_start_address_EN =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h0 ||
	     WILL_FIRE_RL_send_request &&
	     rg_start_address_0_ULT_rg_end_address_4___d35 ;

  // register rg_total_count
  assign rg_total_count_D_IN =
	     MUX_rg_total_count_write_1__SEL_1 ?
	       MUX_rg_total_count_write_1__VAL_1 :
	       MUX_rg_total_count_write_1__VAL_2 ;
  assign rg_total_count_EN =
	     WILL_FIRE_RL_configure_registers &&
	     s_xactor_f_wr_addr_D_OUT[8:5] == 4'h8 ||
	     WILL_FIRE_RL_receive_response ;

  // register rg_word_count
  assign rg_word_count_D_IN = 1'b0 ;
  assign rg_word_count_EN = 1'b0 ;

  // submodule ff_lower_order_bits
  assign ff_lower_order_bits_D_IN = rg_start_address[2:0] ;
  assign ff_lower_order_bits_ENQ = MUX_rg_start_address_write_1__SEL_2 ;
  assign ff_lower_order_bits_DEQ = CAN_FIRE_RL_receive_response ;
  assign ff_lower_order_bits_CLR = 1'b0 ;

  // submodule m_xactor_f_rd_addr
  assign m_xactor_f_rd_addr_D_IN = { rg_start_address, 5'd6 } ;
  assign m_xactor_f_rd_addr_ENQ = MUX_rg_start_address_write_1__SEL_2 ;
  assign m_xactor_f_rd_addr_DEQ =
	     m_xactor_f_rd_addr_EMPTY_N && master_m_arready_arready ;
  assign m_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule m_xactor_f_rd_data
  assign m_xactor_f_rd_data_D_IN =
	     { master_m_rvalid_rresp, master_m_rvalid_rdata } ;
  assign m_xactor_f_rd_data_ENQ =
	     master_m_rvalid_rvalid && m_xactor_f_rd_data_FULL_N ;
  assign m_xactor_f_rd_data_DEQ = CAN_FIRE_RL_receive_response ;
  assign m_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule m_xactor_f_wr_addr
  assign m_xactor_f_wr_addr_D_IN = 37'h0 ;
  assign m_xactor_f_wr_addr_ENQ = 1'b0 ;
  assign m_xactor_f_wr_addr_DEQ =
	     m_xactor_f_wr_addr_EMPTY_N && master_m_awready_awready ;
  assign m_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule m_xactor_f_wr_data
  assign m_xactor_f_wr_data_D_IN = 72'h0 ;
  assign m_xactor_f_wr_data_ENQ = 1'b0 ;
  assign m_xactor_f_wr_data_DEQ =
	     m_xactor_f_wr_data_EMPTY_N && master_m_wready_wready ;
  assign m_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule m_xactor_f_wr_resp
  assign m_xactor_f_wr_resp_D_IN = master_m_bvalid_bresp ;
  assign m_xactor_f_wr_resp_ENQ =
	     master_m_bvalid_bvalid && m_xactor_f_wr_resp_FULL_N ;
  assign m_xactor_f_wr_resp_DEQ = 1'b0 ;
  assign m_xactor_f_wr_resp_CLR = 1'b0 ;

  // submodule s_xactor_f_rd_addr
  assign s_xactor_f_rd_addr_D_IN =
	     { slave_m_arvalid_araddr,
	       slave_m_arvalid_arprot,
	       slave_m_arvalid_arsize } ;
  assign s_xactor_f_rd_addr_ENQ =
	     slave_m_arvalid_arvalid && s_xactor_f_rd_addr_FULL_N ;
  assign s_xactor_f_rd_addr_DEQ = 1'b0 ;
  assign s_xactor_f_rd_addr_CLR = 1'b0 ;

  // submodule s_xactor_f_rd_data
  assign s_xactor_f_rd_data_D_IN = 66'h0 ;
  assign s_xactor_f_rd_data_ENQ = 1'b0 ;
  assign s_xactor_f_rd_data_DEQ =
	     slave_m_rready_rready && s_xactor_f_rd_data_EMPTY_N ;
  assign s_xactor_f_rd_data_CLR = 1'b0 ;

  // submodule s_xactor_f_wr_addr
  assign s_xactor_f_wr_addr_D_IN =
	     { slave_m_awvalid_awaddr,
	       slave_m_awvalid_awprot,
	       slave_m_awvalid_awsize } ;
  assign s_xactor_f_wr_addr_ENQ =
	     slave_m_awvalid_awvalid && s_xactor_f_wr_addr_FULL_N ;
  assign s_xactor_f_wr_addr_DEQ = CAN_FIRE_RL_configure_registers ;
  assign s_xactor_f_wr_addr_CLR = 1'b0 ;

  // submodule s_xactor_f_wr_data
  assign s_xactor_f_wr_data_D_IN =
	     { slave_m_wvalid_wdata, slave_m_wvalid_wstrb } ;
  assign s_xactor_f_wr_data_ENQ =
	     slave_m_wvalid_wvalid && s_xactor_f_wr_data_FULL_N ;
  assign s_xactor_f_wr_data_DEQ = CAN_FIRE_RL_configure_registers ;
  assign s_xactor_f_wr_data_CLR = 1'b0 ;

  // submodule s_xactor_f_wr_resp
  always@(s_xactor_f_wr_addr_D_OUT)
  begin
    case (s_xactor_f_wr_addr_D_OUT[8:5])
      4'h0, 4'h8: s_xactor_f_wr_resp_D_IN = 2'd0;
      default: s_xactor_f_wr_resp_D_IN = 2'd2;
    endcase
  end
  assign s_xactor_f_wr_resp_ENQ = CAN_FIRE_RL_configure_registers ;
  assign s_xactor_f_wr_resp_DEQ =
	     slave_m_bready_bready && s_xactor_f_wr_resp_EMPTY_N ;
  assign s_xactor_f_wr_resp_CLR = 1'b0 ;

  // remaining internal signals
  assign lv_shift__h2655 = { ff_lower_order_bits_D_OUT, 3'd0 } ;
  assign m_xactor_f_rd_dataD_OUT_BITS_63_TO_0_SRL_lv_s_ETC__q2 =
	     m_xactor_f_rd_data_D_OUT[63:0] >> lv_shift__h2655 ;
  assign rg_cnt_ULT_5___d2 = rg_cnt < 5'd5 ;
  assign rg_start_address_0_ULT_rg_end_address_4___d35 =
	     rg_start_address < rg_end_address ;
  assign s_xactor_f_wr_dataD_OUT_BITS_39_TO_8_MINUS_rg_ETC__q1 =
	     s_xactor_f_wr_data_D_OUT[39:8] - rg_start_address ;

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        dataarray_0 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	dataarray_1 <= `BSV_ASSIGNMENT_DELAY 32'd0;
	dump <= `BSV_ASSIGNMENT_DELAY 32'd0;
	rg_cnt <= `BSV_ASSIGNMENT_DELAY 5'd0;
	rg_end_address <= `BSV_ASSIGNMENT_DELAY 32'd0;
	rg_end_sim <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_start <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_start_address <= `BSV_ASSIGNMENT_DELAY 32'd0;
	rg_total_count <= `BSV_ASSIGNMENT_DELAY 32'd0;
	rg_word_count <= `BSV_ASSIGNMENT_DELAY 1'd1;
      end
    else
      begin
        if (dataarray_0_EN)
	  dataarray_0 <= `BSV_ASSIGNMENT_DELAY dataarray_0_D_IN;
	if (dataarray_1_EN)
	  dataarray_1 <= `BSV_ASSIGNMENT_DELAY dataarray_1_D_IN;
	if (dump_EN) dump <= `BSV_ASSIGNMENT_DELAY dump_D_IN;
	if (rg_cnt_EN) rg_cnt <= `BSV_ASSIGNMENT_DELAY rg_cnt_D_IN;
	if (rg_end_address_EN)
	  rg_end_address <= `BSV_ASSIGNMENT_DELAY rg_end_address_D_IN;
	if (rg_end_sim_EN)
	  rg_end_sim <= `BSV_ASSIGNMENT_DELAY rg_end_sim_D_IN;
	if (rg_start_EN) rg_start <= `BSV_ASSIGNMENT_DELAY rg_start_D_IN;
	if (rg_start_address_EN)
	  rg_start_address <= `BSV_ASSIGNMENT_DELAY rg_start_address_D_IN;
	if (rg_total_count_EN)
	  rg_total_count <= `BSV_ASSIGNMENT_DELAY rg_total_count_D_IN;
	if (rg_word_count_EN)
	  rg_word_count <= `BSV_ASSIGNMENT_DELAY rg_word_count_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    dataarray_0 = 32'hAAAAAAAA;
    dataarray_1 = 32'hAAAAAAAA;
    dump = 32'hAAAAAAAA;
    rg_cnt = 5'h0A;
    rg_end_address = 32'hAAAAAAAA;
    rg_end_sim = 1'h0;
    rg_start = 1'h0;
    rg_start_address = 32'hAAAAAAAA;
    rg_total_count = 32'hAAAAAAAA;
    rg_word_count = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_open_file)
	begin
	  TASK_fopen___d3 = $fopen("signature", "w");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_open_file && TASK_fopen___d3 == 32'd0)
	$display("cannot open %s", "signature");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_open_file && TASK_fopen___d3 == 32'd0) $finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_receive_response)
	$fwrite(dump,
		"%4h\n",
		m_xactor_f_rd_dataD_OUT_BITS_63_TO_0_SRL_lv_s_ETC__q2[31:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_receive_response &&
	  m_xactor_f_rd_data_D_OUT[65:64] != 2'd0)
	begin
	  v__h2897 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_receive_response &&
	  m_xactor_f_rd_data_D_OUT[65:64] != 2'd0)
	$display(v__h2897, "\tSIGNATUREDUMP got Bus Error");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_receive_response &&
	  m_xactor_f_rd_data_D_OUT[65:64] != 2'd0)
	$finish(32'd0);
  end
  // synopsys translate_on
endmodule  // mksign_dump_axi4lite

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:06 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// inst_request_get               O    66
// RDY_inst_request_get           O     1
// RDY_inst_response_put          O     1 reg
// tx_stage1_operands_enq_ena     O     1
// tx_stage1_operands_enq_data    O   128
// tx_stage1_meta_enq_ena         O     1
// tx_stage1_meta_enq_data        O    65
// tx_stage1_control_enq_ena      O     1
// tx_stage1_control_enq_data     O    66 reg
// tx_stage1_dump_enq_ena         O     1
// tx_stage1_dump_enq_data        O    96
// RDY_commit_rd_put              O     1
// RDY_ma_update_eEpoch           O     1 const
// RDY_ma_update_wEpoch           O     1 const
// resetpc                        I    64
// CLK                            I     1 clock
// RST_N                          I     1 reset
// inst_response_put              I    35 reg
// tx_stage1_operands_notFull_b   I     1 unused
// tx_stage1_operands_enq_rdy_b   I     1
// tx_stage1_meta_notFull_b       I     1 unused
// tx_stage1_meta_enq_rdy_b       I     1
// tx_stage1_control_notFull_b    I     1 unused
// tx_stage1_control_enq_rdy_b    I     1
// tx_stage1_dump_notFull_b       I     1 unused
// tx_stage1_dump_enq_rdy_b       I     1
// commit_rd_put                  I    69
// ma_flush_newpc                 I    64
// ma_csr_misa_c_c                I     1
// ma_interrupt_i                 I     1
// ma_csr_decode_c                I   152
// ma_trigger_data1_t             I    44
// ma_trigger_data2_t             I   128
// ma_trigger_enable_t            I     2
// EN_inst_response_put           I     1
// EN_commit_rd_put               I     1
// EN_ma_flush                    I     1
// EN_ma_update_eEpoch            I     1
// EN_ma_update_wEpoch            I     1
// EN_inst_request_get            I     1
//
// Combinational paths from inputs to outputs:
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_operands_enq_ena
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    commit_rd_put,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_commit_rd_put,
//    EN_ma_flush) -> tx_stage1_operands_enq_data
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_meta_enq_ena
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    ma_trigger_data1_t,
//    ma_trigger_data2_t,
//    ma_trigger_enable_t,
//    EN_ma_flush) -> tx_stage1_meta_enq_data
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_control_enq_ena
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_control_enq_data
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_dump_enq_ena
//   (tx_stage1_operands_enq_rdy_b,
//    tx_stage1_meta_enq_rdy_b,
//    tx_stage1_control_enq_rdy_b,
//    tx_stage1_dump_enq_rdy_b,
//    ma_csr_misa_c_c,
//    ma_csr_decode_c,
//    EN_ma_flush) -> tx_stage1_dump_enq_data
//
//
// module: This Module implements the instruction-fetch + decode + operand-fetch   functionality of the pipeline.     1. Instruction-Fetch phase:  It generates the new PC, sends the PC to the fabric and in   return expects the instruction response from the fabric. The PC is updated  either when a flush is received from any of the later stages or is simple incremented by 4 or 2  (in case of compressed instructions)    2. Decode phase: Once the instruction is received, it is checked if the instruction is a  compressed instruction or not. If so, then it passes through a decompressor which then converts  the compressed instruction into its 32-bit equivalent encoding. The 32-bit instructions are  then decoded to capture various informations. Most of the decoded information which holds  control-flow information is passed on to the next stage for execution.    3. Operand Fetch: The operand addresses are generated by the decoder and then used to access the  register file. The registerfile itself forward the data of the commit happening in the same  cycle. The fetched operands are then passed on to the next stage.    4. The debugger also is given access to the registerfile through this module.    5. Triggers are also supported to capture events related to program counter or instruction match
//
// Comments on the inlined module `v_trigger_enable':
//   vector: Array of wires capturing which triggers are enabled currently
//
// Comments on the inlined module `v_trigger_data2':
//   vector: Array of wires capturing the tdata2 values from csr
//
// Comments on the inlined module `v_trigger_data1':
//   vector: Array of wires capturing the tdata1 values from csr
//
// Comments on the inlined module `integer_rf':
//   submod: operand register file
//
// Comments on the inlined module `wr_interrupt':
//   wire: This wire will be set if any interrupts have been detected by the core
//
// Comments on the inlined module `wr_csr_decode':
//   wire: this wire caries the current value of certain csrs
//
// Comments on the inlined module `wr_csr_misa_c':
//   wire: this wire carries the current value of the misa_c csr field
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkstage1(resetpc,
		CLK,
		RST_N,

		EN_inst_request_get,
		inst_request_get,
		RDY_inst_request_get,

		inst_response_put,
		EN_inst_response_put,
		RDY_inst_response_put,

		tx_stage1_operands_notFull_b,

		tx_stage1_operands_enq_rdy_b,

		tx_stage1_operands_enq_ena,

		tx_stage1_operands_enq_data,

		tx_stage1_meta_notFull_b,

		tx_stage1_meta_enq_rdy_b,

		tx_stage1_meta_enq_ena,

		tx_stage1_meta_enq_data,

		tx_stage1_control_notFull_b,

		tx_stage1_control_enq_rdy_b,

		tx_stage1_control_enq_ena,

		tx_stage1_control_enq_data,

		tx_stage1_dump_notFull_b,

		tx_stage1_dump_enq_rdy_b,

		tx_stage1_dump_enq_ena,

		tx_stage1_dump_enq_data,

		commit_rd_put,
		EN_commit_rd_put,
		RDY_commit_rd_put,

		ma_flush_newpc,
		EN_ma_flush,

		ma_csr_misa_c_c,

		ma_interrupt_i,

		ma_csr_decode_c,

		EN_ma_update_eEpoch,
		RDY_ma_update_eEpoch,

		EN_ma_update_wEpoch,
		RDY_ma_update_wEpoch,

		ma_trigger_data1_t,

		ma_trigger_data2_t,

		ma_trigger_enable_t);
  input  [63 : 0] resetpc;
  input  CLK;
  input  RST_N;

  // actionvalue method inst_request_get
  input  EN_inst_request_get;
  output [65 : 0] inst_request_get;
  output RDY_inst_request_get;

  // action method inst_response_put
  input  [34 : 0] inst_response_put;
  input  EN_inst_response_put;
  output RDY_inst_response_put;

  // action method tx_stage1_operands_notFull
  input  tx_stage1_operands_notFull_b;

  // action method tx_stage1_operands_enq_rdy
  input  tx_stage1_operands_enq_rdy_b;

  // value method tx_stage1_operands_enq_ena
  output tx_stage1_operands_enq_ena;

  // value method tx_stage1_operands_enq_data
  output [127 : 0] tx_stage1_operands_enq_data;

  // action method tx_stage1_meta_notFull
  input  tx_stage1_meta_notFull_b;

  // action method tx_stage1_meta_enq_rdy
  input  tx_stage1_meta_enq_rdy_b;

  // value method tx_stage1_meta_enq_ena
  output tx_stage1_meta_enq_ena;

  // value method tx_stage1_meta_enq_data
  output [64 : 0] tx_stage1_meta_enq_data;

  // action method tx_stage1_control_notFull
  input  tx_stage1_control_notFull_b;

  // action method tx_stage1_control_enq_rdy
  input  tx_stage1_control_enq_rdy_b;

  // value method tx_stage1_control_enq_ena
  output tx_stage1_control_enq_ena;

  // value method tx_stage1_control_enq_data
  output [65 : 0] tx_stage1_control_enq_data;

  // action method tx_stage1_dump_notFull
  input  tx_stage1_dump_notFull_b;

  // action method tx_stage1_dump_enq_rdy
  input  tx_stage1_dump_enq_rdy_b;

  // value method tx_stage1_dump_enq_ena
  output tx_stage1_dump_enq_ena;

  // value method tx_stage1_dump_enq_data
  output [95 : 0] tx_stage1_dump_enq_data;

  // action method commit_rd_put
  input  [68 : 0] commit_rd_put;
  input  EN_commit_rd_put;
  output RDY_commit_rd_put;

  // action method ma_flush
  input  [63 : 0] ma_flush_newpc;
  input  EN_ma_flush;

  // action method ma_csr_misa_c
  input  ma_csr_misa_c_c;

  // action method ma_interrupt
  input  ma_interrupt_i;

  // action method ma_csr_decode
  input  [151 : 0] ma_csr_decode_c;

  // action method ma_update_eEpoch
  input  EN_ma_update_eEpoch;
  output RDY_ma_update_eEpoch;

  // action method ma_update_wEpoch
  input  EN_ma_update_wEpoch;
  output RDY_ma_update_wEpoch;

  // action method ma_trigger_data1
  input  [43 : 0] ma_trigger_data1_t;

  // action method ma_trigger_data2
  input  [127 : 0] ma_trigger_data2_t;

  // action method ma_trigger_enable
  input  [1 : 0] ma_trigger_enable_t;

  // signals for module outputs
  wire [127 : 0] tx_stage1_operands_enq_data;
  wire [95 : 0] tx_stage1_dump_enq_data;
  wire [65 : 0] inst_request_get, tx_stage1_control_enq_data;
  wire [64 : 0] tx_stage1_meta_enq_data;
  wire RDY_commit_rd_put,
       RDY_inst_request_get,
       RDY_inst_response_put,
       RDY_ma_update_eEpoch,
       RDY_ma_update_wEpoch,
       tx_stage1_control_enq_ena,
       tx_stage1_dump_enq_ena,
       tx_stage1_meta_enq_ena,
       tx_stage1_operands_enq_ena;

  // inlined wires
  reg [21 : 0] v_trigger_data1_0_wget, v_trigger_data1_1_wget;
  wire [151 : 0] wr_csr_decode_wget;
  wire [64 : 0] ff_stage1_meta_w_data_wget;
  wire [63 : 0] rg_fabric_request_port0__write_1,
		rg_fabric_request_port1__read,
		rg_fabric_request_port1__write_1,
		rg_fabric_request_port2__read;
  wire integer_rf_wr_write_address_whas,
       integer_rf_wr_write_data_whas,
       rg_fabric_request_EN_port1__write;

  // register rg_action
  // reg: This register implements a simple state - machine which indicates how the     instruction should be extracted from the cache response.
  reg rg_action;
  wire rg_action_D_IN, rg_action_EN;

  // register rg_discard_lower
  reg rg_discard_lower;
  wire rg_discard_lower_D_IN, rg_discard_lower_EN;

  // register rg_eEpoch
  // reg: holds the current epoch values controlled by the stage2.
  reg rg_eEpoch;
  wire rg_eEpoch_D_IN, rg_eEpoch_EN;

  // register rg_fabric_request
  // reg: register to hold the address of the next request to the fabric.
  reg [63 : 0] rg_fabric_request;
  wire [63 : 0] rg_fabric_request_D_IN;
  wire rg_fabric_request_EN;

  // register rg_index
  // reg: index into the Regfile during initialization sequence.
  reg [4 : 0] rg_index;
  wire [4 : 0] rg_index_D_IN;
  wire rg_index_EN;

  // register rg_initialize
  // reg: register to indicate that the RegFile is being initialized to all zeros
  reg rg_initialize;
  wire rg_initialize_D_IN, rg_initialize_EN;

  // register rg_pc
  // reg: register to hold the PC value of the instruction to be decoded.
  reg [63 : 0] rg_pc;
  reg [63 : 0] rg_pc_D_IN;
  wire rg_pc_EN;

  // register rg_prev
  reg [17 : 0] rg_prev;
  wire [17 : 0] rg_prev_D_IN;
  wire rg_prev_EN;

  // register rg_wEpoch
  // reg: holds the current epoch values controlled by the stage3.
  reg rg_wEpoch;
  wire rg_wEpoch_D_IN, rg_wEpoch_EN;

  // register rg_wfi
  // reg: this is register it set to True when a WFI instruction is executed. It set to     False, when an interrupt has been received or there is a flush from the write - back stage.
  reg rg_wfi;
  wire rg_wfi_D_IN, rg_wfi_EN;

  // ports of submodule ff_memory_response
  wire [34 : 0] ff_memory_response_D_IN, ff_memory_response_D_OUT;
  wire ff_memory_response_CLR,
       ff_memory_response_DEQ,
       ff_memory_response_EMPTY_N,
       ff_memory_response_ENQ,
       ff_memory_response_FULL_N;

  // ports of submodule integer_rf_rf
  wire [63 : 0] integer_rf_rf_D_IN,
		integer_rf_rf_D_OUT_1,
		integer_rf_rf_D_OUT_2;
  wire [4 : 0] integer_rf_rf_ADDR_1,
	       integer_rf_rf_ADDR_2,
	       integer_rf_rf_ADDR_3,
	       integer_rf_rf_ADDR_4,
	       integer_rf_rf_ADDR_5,
	       integer_rf_rf_ADDR_IN;
  wire integer_rf_rf_WE;

  // rule scheduling signals
  wire CAN_FIRE_RL_initialize_regfile,
       CAN_FIRE_RL_process_instruction,
       CAN_FIRE_RL_wait_for_interrupt,
       CAN_FIRE_commit_rd_put,
       CAN_FIRE_inst_request_get,
       CAN_FIRE_inst_response_put,
       CAN_FIRE_ma_csr_decode,
       CAN_FIRE_ma_csr_misa_c,
       CAN_FIRE_ma_flush,
       CAN_FIRE_ma_interrupt,
       CAN_FIRE_ma_trigger_data1,
       CAN_FIRE_ma_trigger_data2,
       CAN_FIRE_ma_trigger_enable,
       CAN_FIRE_ma_update_eEpoch,
       CAN_FIRE_ma_update_wEpoch,
       CAN_FIRE_tx_stage1_control_enq_rdy,
       CAN_FIRE_tx_stage1_control_notFull,
       CAN_FIRE_tx_stage1_dump_enq_rdy,
       CAN_FIRE_tx_stage1_dump_notFull,
       CAN_FIRE_tx_stage1_meta_enq_rdy,
       CAN_FIRE_tx_stage1_meta_notFull,
       CAN_FIRE_tx_stage1_operands_enq_rdy,
       CAN_FIRE_tx_stage1_operands_notFull,
       WILL_FIRE_RL_initialize_regfile,
       WILL_FIRE_RL_process_instruction,
       WILL_FIRE_RL_wait_for_interrupt,
       WILL_FIRE_commit_rd_put,
       WILL_FIRE_inst_request_get,
       WILL_FIRE_inst_response_put,
       WILL_FIRE_ma_csr_decode,
       WILL_FIRE_ma_csr_misa_c,
       WILL_FIRE_ma_flush,
       WILL_FIRE_ma_interrupt,
       WILL_FIRE_ma_trigger_data1,
       WILL_FIRE_ma_trigger_data2,
       WILL_FIRE_ma_trigger_enable,
       WILL_FIRE_ma_update_eEpoch,
       WILL_FIRE_ma_update_wEpoch,
       WILL_FIRE_tx_stage1_control_enq_rdy,
       WILL_FIRE_tx_stage1_control_notFull,
       WILL_FIRE_tx_stage1_dump_enq_rdy,
       WILL_FIRE_tx_stage1_dump_notFull,
       WILL_FIRE_tx_stage1_meta_enq_rdy,
       WILL_FIRE_tx_stage1_meta_notFull,
       WILL_FIRE_tx_stage1_operands_enq_rdy,
       WILL_FIRE_tx_stage1_operands_notFull;

  // inputs to muxes for submodule ports
  wire [63 : 0] MUX_rg_fabric_request_port1__write_1__VAL_2,
		MUX_rg_pc_write_1__VAL_1;
  wire MUX_rg_discard_lower_write_1__SEL_1,
       MUX_rg_fabric_request_port1__write_1__SEL_1,
       MUX_rg_pc_write_1__SEL_1,
       MUX_rg_wfi_write_1__SEL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d446;
  reg TASK_testplusargs___d447;
  reg TASK_testplusargs___d448;
  reg [63 : 0] v__h8601;
  reg TASK_testplusargs___d459;
  reg TASK_testplusargs___d460;
  reg TASK_testplusargs___d461;
  reg [63 : 0] v__h8998;
  reg TASK_testplusargs___d2;
  reg TASK_testplusargs___d3;
  reg TASK_testplusargs___d4;
  reg [63 : 0] v__h2955;
  reg TASK_testplusargs___d17;
  reg TASK_testplusargs___d18;
  reg TASK_testplusargs___d19;
  reg [63 : 0] v__h3340;
  reg TASK_testplusargs___d91;
  reg TASK_testplusargs___d92;
  reg TASK_testplusargs___d93;
  reg [63 : 0] v__h3536;
  reg TASK_testplusargs___d108;
  reg TASK_testplusargs___d109;
  reg TASK_testplusargs___d110;
  reg [63 : 0] v__h4359;
  reg TASK_testplusargs___d116;
  reg TASK_testplusargs___d117;
  reg TASK_testplusargs___d118;
  reg [63 : 0] v__h4531;
  reg TASK_testplusargs___d168;
  reg TASK_testplusargs___d169;
  reg TASK_testplusargs___d170;
  reg [63 : 0] v__h5120;
  reg TASK_testplusargs___d205;
  reg TASK_testplusargs___d206;
  reg TASK_testplusargs___d207;
  reg [63 : 0] v__h5546;
  reg TASK_testplusargs___d212;
  reg TASK_testplusargs___d213;
  reg TASK_testplusargs___d214;
  reg [63 : 0] v__h5785;
  reg TASK_testplusargs___d222;
  reg TASK_testplusargs___d223;
  reg TASK_testplusargs___d224;
  reg [63 : 0] v__h6064;
  reg TASK_testplusargs___d259;
  reg TASK_testplusargs___d260;
  reg TASK_testplusargs___d261;
  reg [63 : 0] v__h6412;
  reg TASK_testplusargs___d266;
  reg TASK_testplusargs___d267;
  reg TASK_testplusargs___d268;
  reg [63 : 0] v__h6581;
  reg TASK_testplusargs___d388;
  reg TASK_testplusargs___d389;
  reg TASK_testplusargs___d390;
  reg [63 : 0] v__h7686;
  reg TASK_testplusargs___d395;
  reg TASK_testplusargs___d396;
  reg TASK_testplusargs___d397;
  reg [63 : 0] v__h7835;
  reg NOT_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_mem_ETC___d96;
  reg TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d114;
  reg TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d115;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194;
  reg TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195;
  reg TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d219;
  reg TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d221;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248;
  reg TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249;
  reg TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d273;
  reg TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d275;
  reg NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393;
  reg NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d400;
  // synopsys translate_on

  // remaining internal signals
  reg [1 : 0] CASE_IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ETC__q5,
	      CASE_decoder_func_32_58_BITS_42_TO_41_0_decode_ETC__q4,
	      IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425;
  reg CASE_v_trigger_data1_0wget_BITS_14_TO_11_2_IF_ETC__q2,
      IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327,
      IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352,
      IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355;
  wire [64 : 0] decoder_func_32___d158;
  wire [63 : 0] _theResult____h6904,
		_theResult____h7088,
		compare_value__h6967,
		ma_trigger_data2_t_BITS_127_TO_64__q3,
		ma_trigger_data2_t_BITS_63_TO_0__q1,
		trigger_compare__h6903,
		trigger_compare__h7087,
		x__h6807,
		x__h7258,
		x__read__h1087,
		x_wget__h1076;
  wire [45 : 0] IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d376;
  wire [31 : 0] _theResult_____4__h4464,
		decode_instruction___1__h4590,
		final_instruction___1__h4584,
		final_instruction__h4155,
		y_avValue_snd_fst__h4179,
		y_avValue_snd_fst__h4187,
		y_avValue_snd_fst__h4189,
		y_avValue_snd_fst__h4209,
		y_avValue_snd_fst__h4211,
		y_avValue_snd_fst__h4240,
		y_avValue_snd_fst__h4244;
  wire [15 : 0] x1_avValue_snd_snd_instruction__h4207,
		x1_avValue_snd_snd_instruction__h4252,
		x1_avValue_snd_snd_instruction__h4254,
		x1_avValue_snd_snd_snd_instruction__h4235,
		x1_avValue_snd_snd_snd_instruction__h4256,
		x1_avValue_snd_snd_snd_instruction__h4258,
		x_instruction__h4177;
  wire [11 : 0] x__h4889;
  wire [7 : 0] chk_interrupt___d152;
  wire [6 : 0] _theResult_____2_meta_funct__h7358,
	       _theResult___fst__h4906,
	       func_cause___1__h4899,
	       x1_avValue_meta_funct__h4765;
  wire [4 : 0] x__read__h1016, x_wget__h1005;
  wire [3 : 0] IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d358;
  wire [1 : 0] IF_wr_csr_decode_wget__41_BITS_151_TO_150_42_E_ETC___d144,
	       curr_epoch__h2865;
  wire IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124,
       IF_chk_interrupt_52_BIT_1_53_OR_ff_memory_resp_ETC___d167,
       IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311,
       IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348,
       IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306,
       IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d326,
       IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340,
       IF_v_trigger_enable_1_wget__72_AND_v_trigger_d_ETC___d356,
       NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277,
       NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d383,
       NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d165,
       NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d86,
       NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d316,
       NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318,
       NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d330,
       NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350,
       decode_word32___d374,
       ff_memory_response_i_notEmpty__3_AND_wr_csr_de_ETC___d47,
       rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65,
       rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d90,
       rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59,
       v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346;

  // actionvalue method inst_request_get
  assign inst_request_get = { rg_fabric_request, curr_epoch__h2865 } ;
  assign RDY_inst_request_get = !rg_initialize ;
  assign CAN_FIRE_inst_request_get = !rg_initialize ;
  assign WILL_FIRE_inst_request_get = EN_inst_request_get ;

  // action method inst_response_put
  assign RDY_inst_response_put = ff_memory_response_FULL_N ;
  assign CAN_FIRE_inst_response_put = ff_memory_response_FULL_N ;
  assign WILL_FIRE_inst_response_put = EN_inst_response_put ;

  // action method tx_stage1_operands_notFull
  assign CAN_FIRE_tx_stage1_operands_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage1_operands_notFull = 1'd1 ;

  // action method tx_stage1_operands_enq_rdy
  assign CAN_FIRE_tx_stage1_operands_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage1_operands_enq_rdy = 1'd1 ;

  // value method tx_stage1_operands_enq_ena
  assign tx_stage1_operands_enq_ena = MUX_rg_pc_write_1__SEL_1 ;

  // value method tx_stage1_operands_enq_data
  assign tx_stage1_operands_enq_data = { x__h6807, x__h7258 } ;

  // action method tx_stage1_meta_notFull
  assign CAN_FIRE_tx_stage1_meta_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage1_meta_notFull = 1'd1 ;

  // action method tx_stage1_meta_enq_rdy
  assign CAN_FIRE_tx_stage1_meta_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage1_meta_enq_rdy = 1'd1 ;

  // value method tx_stage1_meta_enq_ena
  assign tx_stage1_meta_enq_ena = MUX_rg_pc_write_1__SEL_1 ;

  // value method tx_stage1_meta_enq_data
  assign tx_stage1_meta_enq_data =
	     { ff_stage1_meta_w_data_wget[64:43],
	       CASE_IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ETC__q5,
	       ff_stage1_meta_w_data_wget[40:0] } ;

  // action method tx_stage1_control_notFull
  assign CAN_FIRE_tx_stage1_control_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage1_control_notFull = 1'd1 ;

  // action method tx_stage1_control_enq_rdy
  assign CAN_FIRE_tx_stage1_control_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage1_control_enq_rdy = 1'd1 ;

  // value method tx_stage1_control_enq_ena
  assign tx_stage1_control_enq_ena = MUX_rg_pc_write_1__SEL_1 ;

  // value method tx_stage1_control_enq_data
  assign tx_stage1_control_enq_data = { curr_epoch__h2865, rg_pc } ;

  // action method tx_stage1_dump_notFull
  assign CAN_FIRE_tx_stage1_dump_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage1_dump_notFull = 1'd1 ;

  // action method tx_stage1_dump_enq_rdy
  assign CAN_FIRE_tx_stage1_dump_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage1_dump_enq_rdy = 1'd1 ;

  // value method tx_stage1_dump_enq_ena
  assign tx_stage1_dump_enq_ena = MUX_rg_pc_write_1__SEL_1 ;

  // value method tx_stage1_dump_enq_data
  assign tx_stage1_dump_enq_data = { rg_pc, final_instruction__h4155 } ;

  // action method commit_rd_put
  assign RDY_commit_rd_put = !rg_initialize ;
  assign CAN_FIRE_commit_rd_put = !rg_initialize ;
  assign WILL_FIRE_commit_rd_put = EN_commit_rd_put ;

  // action method ma_flush
  assign CAN_FIRE_ma_flush = 1'd1 ;
  assign WILL_FIRE_ma_flush = EN_ma_flush ;

  // action method ma_csr_misa_c
  assign CAN_FIRE_ma_csr_misa_c = 1'd1 ;
  assign WILL_FIRE_ma_csr_misa_c = 1'd1 ;

  // action method ma_interrupt
  assign CAN_FIRE_ma_interrupt = 1'd1 ;
  assign WILL_FIRE_ma_interrupt = 1'd1 ;

  // action method ma_csr_decode
  assign CAN_FIRE_ma_csr_decode = 1'd1 ;
  assign WILL_FIRE_ma_csr_decode = 1'd1 ;

  // action method ma_update_eEpoch
  assign RDY_ma_update_eEpoch = 1'd1 ;
  assign CAN_FIRE_ma_update_eEpoch = 1'd1 ;
  assign WILL_FIRE_ma_update_eEpoch = EN_ma_update_eEpoch ;

  // action method ma_update_wEpoch
  assign RDY_ma_update_wEpoch = 1'd1 ;
  assign CAN_FIRE_ma_update_wEpoch = 1'd1 ;
  assign WILL_FIRE_ma_update_wEpoch = EN_ma_update_wEpoch ;

  // action method ma_trigger_data1
  assign CAN_FIRE_ma_trigger_data1 = 1'd1 ;
  assign WILL_FIRE_ma_trigger_data1 = 1'd1 ;

  // action method ma_trigger_data2
  assign CAN_FIRE_ma_trigger_data2 = 1'd1 ;
  assign WILL_FIRE_ma_trigger_data2 = 1'd1 ;

  // action method ma_trigger_enable
  assign CAN_FIRE_ma_trigger_enable = 1'd1 ;
  assign WILL_FIRE_ma_trigger_enable = 1'd1 ;

  // submodule ff_memory_response
  // fifo: to hold the instruction response from the fabric
  FIFO2 #(.width(32'd35), .guarded(32'd1)) ff_memory_response(.RST(RST_N),
							      .CLK(CLK),
							      .D_IN(ff_memory_response_D_IN),
							      .ENQ(ff_memory_response_ENQ),
							      .DEQ(ff_memory_response_DEQ),
							      .CLR(ff_memory_response_CLR),
							      .D_OUT(ff_memory_response_D_OUT),
							      .FULL_N(ff_memory_response_FULL_N),
							      .EMPTY_N(ff_memory_response_EMPTY_N));

  // submodule integer_rf_rf
  RegFile #(.addr_width(32'd5),
	    .data_width(32'd64),
	    .lo(5'd0),
	    .hi(5'd31)) integer_rf_rf(.CLK(CLK),
				      .ADDR_1(integer_rf_rf_ADDR_1),
				      .ADDR_2(integer_rf_rf_ADDR_2),
				      .ADDR_3(integer_rf_rf_ADDR_3),
				      .ADDR_4(integer_rf_rf_ADDR_4),
				      .ADDR_5(integer_rf_rf_ADDR_5),
				      .ADDR_IN(integer_rf_rf_ADDR_IN),
				      .D_IN(integer_rf_rf_D_IN),
				      .WE(integer_rf_rf_WE),
				      .D_OUT_1(integer_rf_rf_D_OUT_1),
				      .D_OUT_2(integer_rf_rf_D_OUT_2),
				      .D_OUT_3(),
				      .D_OUT_4(),
				      .D_OUT_5());

  // rule RL_initialize_regfile
  //   rule: initialize all the registers to 0 on reset
  assign CAN_FIRE_RL_initialize_regfile = rg_initialize ;
  assign WILL_FIRE_RL_initialize_regfile = rg_initialize ;

  // rule RL_wait_for_interrupt
  //   rule:This rule is fired when the core has executed the WFI instruction and waiting     for an intterupt to the core to resume fetch
  assign CAN_FIRE_RL_wait_for_interrupt = rg_wfi && !rg_initialize ;
  assign WILL_FIRE_RL_wait_for_interrupt =
	     CAN_FIRE_RL_wait_for_interrupt && !EN_ma_flush ;

  // rule RL_process_instruction
  //   rule:This rule will receive the instruction from the memory subsystem and decide if     the instruction is compressed or not. The final instruction is then sent to the next stage.    To extract the instruction from the memory response a state machine is implemented.        1. First the epochs are compared and if a mis - match is observed then the response is     dropped without any other changes to the state of the module.    2. if rg_discard is set and compressed is enabled then the lower 16 - bits of the    resposne are discarded and the upper 16 - bits are probed to check if it is a compressed    instruction. If so, then the instruction is sent to the next stage. However is it is not a    compressed instruction it means the upper 16 - bits of the response refer to the lower 16 -    bits of a 32 - bit instruction and thus we will have to wait for the next response from the     cache to form the instruction is send to the next stage. To ensure the concatenation happens     in the next response we set rg_action to ChecPrev and set enque_instruction to False.    3. if rg_action is set to None, then we simply probe the lower 2 - bits to the response to    check if it is compressed. If so then the lower 16 bits form an instruction which is sent to    the next stage, the upper 16 - bits are stored to rg_instruction and rg_action is set to    CheckPrev to ensure that in the next resposne we first probe rg_instruction.    4. if rg_Action if set to CheckPrev then we first probe the lower 2 - bits of the     rg_instruction which leads to two possibilities. Either rg_instruction could hold a    compressed instruction from the previous response, in which case the current memory response    is not dequed and rg_instruction is sent to the next stage. This can happen due to state - 3    mentioned above. The other possibility is that rg_instruction holds the lower 16 - bits of a    32 - bit isntruction, in which case we have concatenate the lower 16 - bits of the response     with rg_instruction and send to the next, and also store the upper 16 - bits of the response     into rg_instruction. rg_Action in this case will remain CheckPrev so that the upper bits of     this repsonse are probed in the next cycle.
  assign CAN_FIRE_RL_process_instruction =
	     ff_memory_response_i_notEmpty__3_AND_wr_csr_de_ETC___d47 &&
	     !rg_wfi &&
	     !rg_initialize ;
  assign WILL_FIRE_RL_process_instruction =
	     CAN_FIRE_RL_process_instruction && !EN_ma_flush ;

  // inputs to muxes for submodule ports
  assign MUX_rg_discard_lower_write_1__SEL_1 =
	     WILL_FIRE_RL_process_instruction &&
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d90 ;
  assign MUX_rg_fabric_request_port1__write_1__SEL_1 =
	     rg_initialize && rg_index == 5'd31 ;
  assign MUX_rg_pc_write_1__SEL_1 =
	     WILL_FIRE_RL_process_instruction &&
	     NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277 ;
  assign MUX_rg_wfi_write_1__SEL_1 =
	     WILL_FIRE_RL_wait_for_interrupt && ma_interrupt_i ;
  assign MUX_rg_fabric_request_port1__write_1__VAL_2 =
	     { ma_flush_newpc[63:2], 2'b0 } ;
  assign MUX_rg_pc_write_1__VAL_1 =
	     rg_pc +
	     ((rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	       IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124 &&
	       NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d383 &&
	       ma_csr_misa_c_c) ?
		64'd2 :
		64'd4) ;

  // inlined wires
  assign wr_csr_decode_wget =
	     { (ma_csr_decode_c[151:150] == 2'd3) ?
		 ma_csr_decode_c[151:150] :
		 2'd0,
	       ma_csr_decode_c[149:0] } ;
  assign integer_rf_wr_write_address_whas =
	     rg_initialize || EN_commit_rd_put ;
  assign integer_rf_wr_write_data_whas = EN_commit_rd_put || rg_initialize ;
  assign ff_stage1_meta_w_data_wget =
	     { decoder_func_32___d158[64:47],
	       IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d376,
	       decoder_func_32___d158[0] } ;
  always@(ma_trigger_data1_t)
  begin
    case (ma_trigger_data1_t[21:20])
      2'd0, 2'd1, 2'd2: v_trigger_data1_0_wget = ma_trigger_data1_t[21:0];
      2'd3:
	  v_trigger_data1_0_wget =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(ma_trigger_data1_t)
  begin
    case (ma_trigger_data1_t[43:42])
      2'd0, 2'd1, 2'd2: v_trigger_data1_1_wget = ma_trigger_data1_t[43:22];
      2'd3:
	  v_trigger_data1_1_wget =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  assign rg_fabric_request_port0__write_1 = rg_fabric_request + 64'd4 ;
  assign rg_fabric_request_port1__read =
	     EN_inst_request_get ?
	       rg_fabric_request_port0__write_1 :
	       rg_fabric_request ;
  assign rg_fabric_request_EN_port1__write =
	     rg_initialize && rg_index == 5'd31 || EN_ma_flush ;
  assign rg_fabric_request_port1__write_1 =
	     MUX_rg_fabric_request_port1__write_1__SEL_1 ?
	       resetpc :
	       MUX_rg_fabric_request_port1__write_1__VAL_2 ;
  assign rg_fabric_request_port2__read =
	     rg_fabric_request_EN_port1__write ?
	       rg_fabric_request_port1__write_1 :
	       rg_fabric_request_port1__read ;

  // register rg_action
  assign rg_action_D_IN =
	     !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 ||
	     !rg_action &&
	     rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 ;
  assign rg_action_EN =
	     WILL_FIRE_RL_process_instruction &&
	     (NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d86 ||
	      !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65) ;

  // register rg_discard_lower
  assign rg_discard_lower_D_IN =
	     !MUX_rg_discard_lower_write_1__SEL_1 &&
	     ma_flush_newpc[1:0] != 2'd0 ;
  assign rg_discard_lower_EN =
	     WILL_FIRE_RL_process_instruction &&
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d90 ||
	     EN_ma_flush ;

  // register rg_eEpoch
  assign rg_eEpoch_D_IN = ~rg_eEpoch ;
  assign rg_eEpoch_EN = EN_ma_update_eEpoch ;

  // register rg_fabric_request
  assign rg_fabric_request_D_IN = rg_fabric_request_port2__read ;
  assign rg_fabric_request_EN = 1'b1 ;

  // register rg_index
  assign rg_index_D_IN = rg_index + 5'd1 ;
  assign rg_index_EN = rg_initialize ;

  // register rg_initialize
  assign rg_initialize_D_IN = 1'd0 ;
  assign rg_initialize_EN = MUX_rg_fabric_request_port1__write_1__SEL_1 ;

  // register rg_pc
  always@(MUX_rg_pc_write_1__SEL_1 or
	  MUX_rg_pc_write_1__VAL_1 or
	  MUX_rg_fabric_request_port1__write_1__SEL_1 or
	  resetpc or EN_ma_flush or ma_flush_newpc)
  case (1'b1)
    MUX_rg_pc_write_1__SEL_1: rg_pc_D_IN = MUX_rg_pc_write_1__VAL_1;
    MUX_rg_fabric_request_port1__write_1__SEL_1: rg_pc_D_IN = resetpc;
    EN_ma_flush: rg_pc_D_IN = ma_flush_newpc;
    default: rg_pc_D_IN = 64'hAAAAAAAAAAAAAAAA /* unspecified value */ ;
  endcase
  assign rg_pc_EN =
	     WILL_FIRE_RL_process_instruction &&
	     NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277 ||
	     rg_initialize && rg_index == 5'd31 ||
	     EN_ma_flush ;

  // register rg_prev
  assign rg_prev_D_IN = { x_instruction__h4177, curr_epoch__h2865 } ;
  assign rg_prev_EN = WILL_FIRE_RL_process_instruction ;

  // register rg_wEpoch
  assign rg_wEpoch_D_IN = ~rg_wEpoch ;
  assign rg_wEpoch_EN = EN_ma_update_wEpoch ;

  // register rg_wfi
  assign rg_wfi_D_IN = !MUX_rg_wfi_write_1__SEL_1 && !EN_ma_flush ;
  assign rg_wfi_EN =
	     WILL_FIRE_RL_wait_for_interrupt && ma_interrupt_i ||
	     WILL_FIRE_RL_process_instruction &&
	     IF_chk_interrupt_52_BIT_1_53_OR_ff_memory_resp_ETC___d167 ||
	     EN_ma_flush ;

  // submodule ff_memory_response
  assign ff_memory_response_D_IN = inst_response_put ;
  assign ff_memory_response_ENQ = EN_inst_response_put ;
  assign ff_memory_response_DEQ =
	     WILL_FIRE_RL_process_instruction &&
	     (rg_prev[3:2] == 2'b11 || rg_action ||
	      !rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 ||
	      !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65) ;
  assign ff_memory_response_CLR = 1'b0 ;

  // submodule integer_rf_rf
  assign integer_rf_rf_ADDR_1 = decoder_func_32___d158[59:55] ;
  assign integer_rf_rf_ADDR_2 = decoder_func_32___d158[64:60] ;
  assign integer_rf_rf_ADDR_3 = 5'h0 ;
  assign integer_rf_rf_ADDR_4 = 5'h0 ;
  assign integer_rf_rf_ADDR_5 = 5'h0 ;
  assign integer_rf_rf_ADDR_IN =
	     rg_initialize ? rg_index : commit_rd_put[68:64] ;
  assign integer_rf_rf_D_IN = rg_initialize ? 64'd0 : commit_rd_put[63:0] ;
  assign integer_rf_rf_WE = integer_rf_wr_write_address_whas ;

  // remaining internal signals
  module_fn_decompress instance_fn_decompress_2(.fn_decompress_inst(final_instruction__h4155[15:0]),
						.fn_decompress(decode_instruction___1__h4590));
  module_chk_interrupt instance_chk_interrupt_1(.chk_interrupt_prv(IF_wr_csr_decode_wget__41_BITS_151_TO_150_42_E_ETC___d144),
						.chk_interrupt_mstatus(wr_csr_decode_wget[63:0]),
						.chk_interrupt_mip({ 2'd0,
								     x__h4889 }),
						.chk_interrupt_mie(wr_csr_decode_wget[137:126]),
						.chk_interrupt_mideleg(wr_csr_decode_wget[125:114]),
						.chk_interrupt_uip(wr_csr_decode_wget[113:102]),
						.chk_interrupt_uie(wr_csr_decode_wget[101:90]),
						.chk_interrupt(chk_interrupt___d152));
  module_decoder_func_32 instance_decoder_func_32_3(.decoder_func_32_inst(_theResult_____4__h4464),
						    .decoder_func_32_csrs({ IF_wr_csr_decode_wget__41_BITS_151_TO_150_42_E_ETC___d144,
									    wr_csr_decode_wget[149:0] }),
						    .decoder_func_32_compressed(rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
										IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124),
						    .decoder_func_32(decoder_func_32___d158));
  module_decode_word32 instance_decode_word32_0(.decode_word32_inst(_theResult_____4__h4464),
						.decode_word32_misa_c(wr_csr_decode_wget[66]),
						.decode_word32(decode_word32___d374));
  assign IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d358 =
	     (IF_v_trigger_enable_1_wget__72_AND_v_trigger_d_ETC___d356 ||
	      chk_interrupt___d152[1] ||
	      ff_memory_response_D_OUT[0]) ?
	       4'd6 :
	       decoder_func_32___d158[46:43] ;
  assign IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d376 =
	     { IF_IF_v_trigger_enable_1_wget__72_AND_v_trigge_ETC___d358,
	       CASE_decoder_func_32_58_BITS_42_TO_41_0_decode_ETC__q4,
	       decoder_func_32___d158[40:9],
	       _theResult_____2_meta_funct__h7358,
	       decode_word32___d374 } ;
  assign IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124 =
	     (!rg_action &&
	      rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59) ?
	       rg_prev[3:2] != 2'b11 :
	       ((rg_discard_lower && ma_csr_misa_c_c) ?
		  ff_memory_response_D_OUT[20:19] != 2'b11 :
		  ff_memory_response_D_OUT[4:3] != 2'b11 && ma_csr_misa_c_c) ;
  assign IF_chk_interrupt_52_BIT_1_53_OR_ff_memory_resp_ETC___d167 =
	     ((chk_interrupt___d152[1] || ff_memory_response_D_OUT[0]) ?
		4'd6 :
		decoder_func_32___d158[46:43]) ==
	     4'd7 &&
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	     NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d165 ;
  assign IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311 =
	     trigger_compare__h6903 == _theResult____h6904 ;
  assign IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348 =
	     trigger_compare__h7087 == _theResult____h7088 ||
	     !v_trigger_data1_0_wget[10] &&
	     v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346 ;
  assign IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306 =
	     _theResult____h6904 < trigger_compare__h6903 ;
  assign IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d326 =
	     IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306 ||
	     ((v_trigger_data1_0_wget[14:11] == 4'd2) ?
		!IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306 :
		v_trigger_data1_0_wget[14:11] == 4'd0 &&
		IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311) ;
  assign IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 =
	     _theResult____h7088 < trigger_compare__h7087 ;
  assign IF_v_trigger_enable_1_wget__72_AND_v_trigger_d_ETC___d356 =
	     (ma_trigger_enable_t[1] &&
	      v_trigger_data1_1_wget[21:20] == 2'd0 &&
	      NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d330) ?
	       IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355 :
	       v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346 ;
  assign IF_wr_csr_decode_wget__41_BITS_151_TO_150_42_E_ETC___d144 =
	     (wr_csr_decode_wget[151:150] == 2'd3) ?
	       wr_csr_decode_wget[151:150] :
	       2'd0 ;
  assign NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277 =
	     ((chk_interrupt___d152[1] || ff_memory_response_D_OUT[0]) ?
		4'd6 :
		decoder_func_32___d158[46:43]) !=
	     4'd7 &&
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	     NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d165 ;
  assign NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d383 =
	     ((chk_interrupt___d152[1] || ff_memory_response_D_OUT[0]) ?
		4'd6 :
		decoder_func_32___d158[46:43]) !=
	     4'd7 &&
	     (!rg_action &&
	      rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 ||
	      !rg_discard_lower ||
	      ff_memory_response_D_OUT[20:19] != 2'b11) ;
  assign NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d165 =
	     !rg_action &&
	     rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 ||
	     !rg_discard_lower ||
	     !ma_csr_misa_c_c ||
	     ff_memory_response_D_OUT[20:19] != 2'b11 ;
  assign NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_5__ETC___d86 =
	     !rg_action &&
	     rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 &&
	     rg_prev[3:2] != 2'b11 ||
	     (rg_action ||
	      !rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59) &&
	     (rg_discard_lower && ma_csr_misa_c_c &&
	      ff_memory_response_D_OUT[20:19] == 2'b11 ||
	      !rg_discard_lower && ff_memory_response_D_OUT[4:3] != 2'b11 &&
	      ma_csr_misa_c_c) ;
  assign NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d316 =
	     !ma_trigger_enable_t[0] ||
	     v_trigger_data1_0_wget[21:20] != 2'd0 ||
	     !v_trigger_data1_0_wget[17] ||
	     CASE_v_trigger_data1_0wget_BITS_14_TO_11_2_IF_ETC__q2 ;
  assign NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318 =
	     !ma_trigger_enable_t[0] ||
	     v_trigger_data1_0_wget[21:20] != 2'd0 ||
	     !v_trigger_data1_0_wget[17] ||
	     !v_trigger_data1_0_wget[10] ;
  assign NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d330 =
	     (NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d316 &&
	      NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318 ||
	      ma_trigger_enable_t[0] &&
	      v_trigger_data1_0_wget[21:20] == 2'd0 &&
	      v_trigger_data1_0_wget[17] &&
	      v_trigger_data1_0_wget[10] &&
	      IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327) &&
	     v_trigger_data1_1_wget[17] ;
  assign NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350 =
	     NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318 &&
	     ((v_trigger_data1_1_wget[14:11] == 4'd0) ?
		IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348 :
		v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346) ;
  assign _theResult_____2_meta_funct__h7358 =
	     IF_v_trigger_enable_1_wget__72_AND_v_trigger_d_ETC___d356 ?
	       7'd3 :
	       x1_avValue_meta_funct__h4765 ;
  assign _theResult_____4__h4464 =
	     (rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	      IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124) ?
	       decode_instruction___1__h4590 :
	       final_instruction__h4155 ;
  assign _theResult____h6904 =
	     v_trigger_data1_0_wget[1] ? compare_value__h6967 : rg_pc ;
  assign _theResult____h7088 =
	     v_trigger_data1_1_wget[1] ? compare_value__h6967 : rg_pc ;
  assign _theResult___fst__h4906 =
	     ff_memory_response_D_OUT[0] ?
	       7'd1 :
	       decoder_func_32___d158[8:2] ;
  assign compare_value__h6967 = { 32'd0, _theResult_____4__h4464 } ;
  assign curr_epoch__h2865 = { rg_eEpoch, rg_wEpoch } ;
  assign ff_memory_response_i_notEmpty__3_AND_wr_csr_de_ETC___d47 =
	     ff_memory_response_EMPTY_N && tx_stage1_operands_enq_rdy_b &&
	     tx_stage1_meta_enq_rdy_b &&
	     tx_stage1_control_enq_rdy_b &&
	     tx_stage1_dump_enq_rdy_b ;
  assign final_instruction___1__h4584 =
	     { 16'd0, ff_memory_response_D_OUT[34:19] } ;
  assign final_instruction__h4155 =
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 ?
	       y_avValue_snd_fst__h4179 :
	       32'd0 ;
  assign func_cause___1__h4899 = { 1'd0, chk_interrupt___d152[7:2] } ;
  assign ma_trigger_data2_t_BITS_127_TO_64__q3 = ma_trigger_data2_t[127:64] ;
  assign ma_trigger_data2_t_BITS_63_TO_0__q1 = ma_trigger_data2_t[63:0] ;
  assign rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 =
	     curr_epoch__h2865 == ff_memory_response_D_OUT[2:1] ;
  assign rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d90 =
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	     (rg_action ||
	      !rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59) &&
	     rg_discard_lower &&
	     ma_csr_misa_c_c ;
  assign rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59 =
	     rg_prev[1:0] == curr_epoch__h2865 ;
  assign trigger_compare__h6903 =
	     (rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	      IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124 &&
	      v_trigger_data1_0_wget[5:2] == 4'd2) ?
	       { 48'd0, ma_trigger_data2_t_BITS_63_TO_0__q1[15:0] } :
	       ma_trigger_data2_t[63:0] ;
  assign trigger_compare__h7087 =
	     (rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	      IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124 &&
	      v_trigger_data1_1_wget[5:2] == 4'd2) ?
	       { 48'd0, ma_trigger_data2_t_BITS_127_TO_64__q3[15:0] } :
	       ma_trigger_data2_t[127:64] ;
  assign v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346 =
	     ma_trigger_enable_t[0] &&
	     v_trigger_data1_0_wget[21:20] == 2'd0 &&
	     v_trigger_data1_0_wget[17] &&
	     IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327 ;
  assign x1_avValue_meta_funct__h4765 =
	     chk_interrupt___d152[1] ?
	       func_cause___1__h4899 :
	       _theResult___fst__h4906 ;
  assign x1_avValue_snd_snd_instruction__h4207 =
	     (rg_prev[3:2] == 2'b11) ?
	       ff_memory_response_D_OUT[34:19] :
	       rg_prev[17:2] ;
  assign x1_avValue_snd_snd_instruction__h4252 =
	     ma_csr_misa_c_c ?
	       ff_memory_response_D_OUT[34:19] :
	       rg_prev[17:2] ;
  assign x1_avValue_snd_snd_instruction__h4254 =
	     (ff_memory_response_D_OUT[4:3] == 2'b11) ?
	       rg_prev[17:2] :
	       x1_avValue_snd_snd_instruction__h4252 ;
  assign x1_avValue_snd_snd_snd_instruction__h4235 =
	     (ff_memory_response_D_OUT[20:19] == 2'b11) ?
	       ff_memory_response_D_OUT[34:19] :
	       rg_prev[17:2] ;
  assign x1_avValue_snd_snd_snd_instruction__h4256 =
	     (rg_discard_lower && ma_csr_misa_c_c) ?
	       x1_avValue_snd_snd_snd_instruction__h4235 :
	       x1_avValue_snd_snd_instruction__h4254 ;
  assign x1_avValue_snd_snd_snd_instruction__h4258 =
	     (!rg_action &&
	      rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59) ?
	       x1_avValue_snd_snd_instruction__h4207 :
	       x1_avValue_snd_snd_snd_instruction__h4256 ;
  assign x__h4889 = wr_csr_decode_wget[149:138] ;
  assign x__h6807 =
	     (decoder_func_32___d158[64:60] == x__read__h1016) ?
	       x__read__h1087 :
	       integer_rf_rf_D_OUT_2 ;
  assign x__h7258 =
	     (decoder_func_32___d158[59:55] == x__read__h1016) ?
	       x__read__h1087 :
	       integer_rf_rf_D_OUT_1 ;
  assign x__read__h1016 =
	     integer_rf_wr_write_address_whas ? x_wget__h1005 : 5'd0 ;
  assign x__read__h1087 =
	     integer_rf_wr_write_data_whas ? x_wget__h1076 : 64'd0 ;
  assign x_instruction__h4177 =
	     rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 ?
	       x1_avValue_snd_snd_snd_instruction__h4258 :
	       rg_prev[17:2] ;
  assign x_wget__h1005 = rg_initialize ? rg_index : commit_rd_put[68:64] ;
  assign x_wget__h1076 = EN_commit_rd_put ? commit_rd_put[63:0] : 64'd0 ;
  assign y_avValue_snd_fst__h4179 =
	     (!rg_action &&
	      rg_prev_1_BITS_1_TO_0_5_EQ_rg_eEpoch_6_CONCAT__ETC___d59) ?
	       y_avValue_snd_fst__h4187 :
	       y_avValue_snd_fst__h4189 ;
  assign y_avValue_snd_fst__h4187 =
	     { (rg_prev[3:2] == 2'b11) ?
		 ff_memory_response_D_OUT[18:3] :
		 16'd0,
	       rg_prev[17:2] } ;
  assign y_avValue_snd_fst__h4189 =
	     (rg_discard_lower && ma_csr_misa_c_c) ?
	       y_avValue_snd_fst__h4209 :
	       y_avValue_snd_fst__h4211 ;
  assign y_avValue_snd_fst__h4209 =
	     (ff_memory_response_D_OUT[20:19] == 2'b11) ?
	       32'd0 :
	       final_instruction___1__h4584 ;
  assign y_avValue_snd_fst__h4211 =
	     (ff_memory_response_D_OUT[4:3] == 2'b11) ?
	       ff_memory_response_D_OUT[34:3] :
	       y_avValue_snd_fst__h4240 ;
  assign y_avValue_snd_fst__h4240 =
	     ma_csr_misa_c_c ? y_avValue_snd_fst__h4244 : 32'd0 ;
  assign y_avValue_snd_fst__h4244 =
	     { 16'd0, ff_memory_response_D_OUT[18:3] } ;
  always@(v_trigger_data1_0_wget or
	  IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311 or
	  IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306)
  begin
    case (v_trigger_data1_0_wget[14:11])
      4'd2:
	  CASE_v_trigger_data1_0wget_BITS_14_TO_11_2_IF_ETC__q2 =
	      IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306;
      4'd3:
	  CASE_v_trigger_data1_0wget_BITS_14_TO_11_2_IF_ETC__q2 =
	      !IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306;
      default: CASE_v_trigger_data1_0wget_BITS_14_TO_11_2_IF_ETC__q2 =
		   v_trigger_data1_0_wget[14:11] != 4'd0 ||
		   !IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311;
    endcase
  end
  always@(v_trigger_data1_0_wget or
	  IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311 or
	  IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306 or
	  IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d326)
  begin
    case (v_trigger_data1_0_wget[14:11])
      4'd2:
	  IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327 =
	      !IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d306;
      4'd3:
	  IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327 =
	      IF_v_trigger_data1_0_wget__75_BIT_1_91_THEN_0__ETC___d326;
      default: IF_v_trigger_data1_0_wget__75_BITS_14_TO_11_01_ETC___d327 =
		   v_trigger_data1_0_wget[14:11] == 4'd0 &&
		   IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d311;
    endcase
  end
  always@(v_trigger_data1_1_wget or
	  v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346 or
	  IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348 or
	  IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 or
	  NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350)
  begin
    case (v_trigger_data1_1_wget[14:11])
      4'd0:
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352 =
	      IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348;
      4'd2:
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352 =
	      !IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 ||
	      NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350;
      default: IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352 =
		   v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346;
    endcase
  end
  always@(v_trigger_data1_1_wget or
	  v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346 or
	  IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348 or
	  IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 or
	  NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350 or
	  NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318 or
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352)
  begin
    case (v_trigger_data1_1_wget[14:11])
      4'd0:
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355 =
	      IF_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memo_ETC___d348;
      4'd2:
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355 =
	      !IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 ||
	      NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d350;
      4'd3:
	  IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355 =
	      IF_v_trigger_data1_1_wget__29_BIT_1_45_THEN_0__ETC___d340 ||
	      NOT_v_trigger_enable_0_wget__18_20_OR_NOT_v_tr_ETC___d318 &&
	      IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d352;
      default: IF_v_trigger_data1_1_wget__29_BITS_14_TO_11_55_ETC___d355 =
		   v_trigger_enable_0_wget__18_AND_v_trigger_data_ETC___d346;
    endcase
  end
  always@(decoder_func_32___d158)
  begin
    case (decoder_func_32___d158[42:41])
      2'd0, 2'd1, 2'd3:
	  CASE_decoder_func_32_58_BITS_42_TO_41_0_decode_ETC__q4 =
	      decoder_func_32___d158[42:41];
      2'd2: CASE_decoder_func_32_58_BITS_42_TO_41_0_decode_ETC__q4 = 2'd2;
    endcase
  end
  always@(ff_stage1_meta_w_data_wget)
  begin
    case (ff_stage1_meta_w_data_wget[42:41])
      2'd0, 2'd1:
	  IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425 =
	      ff_stage1_meta_w_data_wget[42:41];
      2'd2: IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425 = 2'd3;
      2'd3: IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425 = 2'd2;
    endcase
  end
  always@(IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425)
  begin
    case (IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425)
      2'd0, 2'd1:
	  CASE_IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ETC__q5 =
	      IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ff_s_ETC___d425;
      2'd2: CASE_IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ETC__q5 = 2'd3;
      2'd3: CASE_IF_ff_stage1_meta_w_data_whas__10_THEN_IF_ETC__q5 = 2'd2;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_action <= `BSV_ASSIGNMENT_DELAY 1'd1;
	rg_discard_lower <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_eEpoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_fabric_request <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_index <= `BSV_ASSIGNMENT_DELAY 5'd0;
	rg_initialize <= `BSV_ASSIGNMENT_DELAY 1'd1;
	rg_pc <= `BSV_ASSIGNMENT_DELAY 64'd0;
	rg_prev <= `BSV_ASSIGNMENT_DELAY 18'd0;
	rg_wEpoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_wfi <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_action_EN) rg_action <= `BSV_ASSIGNMENT_DELAY rg_action_D_IN;
	if (rg_discard_lower_EN)
	  rg_discard_lower <= `BSV_ASSIGNMENT_DELAY rg_discard_lower_D_IN;
	if (rg_eEpoch_EN) rg_eEpoch <= `BSV_ASSIGNMENT_DELAY rg_eEpoch_D_IN;
	if (rg_fabric_request_EN)
	  rg_fabric_request <= `BSV_ASSIGNMENT_DELAY rg_fabric_request_D_IN;
	if (rg_index_EN) rg_index <= `BSV_ASSIGNMENT_DELAY rg_index_D_IN;
	if (rg_initialize_EN)
	  rg_initialize <= `BSV_ASSIGNMENT_DELAY rg_initialize_D_IN;
	if (rg_pc_EN) rg_pc <= `BSV_ASSIGNMENT_DELAY rg_pc_D_IN;
	if (rg_prev_EN) rg_prev <= `BSV_ASSIGNMENT_DELAY rg_prev_D_IN;
	if (rg_wEpoch_EN) rg_wEpoch <= `BSV_ASSIGNMENT_DELAY rg_wEpoch_D_IN;
	if (rg_wfi_EN) rg_wfi <= `BSV_ASSIGNMENT_DELAY rg_wfi_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_action = 1'h0;
    rg_discard_lower = 1'h0;
    rg_eEpoch = 1'h0;
    rg_fabric_request = 64'hAAAAAAAAAAAAAAAA;
    rg_index = 5'h0A;
    rg_initialize = 1'h0;
    rg_pc = 64'hAAAAAAAAAAAAAAAA;
    rg_prev = 18'h2AAAA;
    rg_wEpoch = 1'h0;
    rg_wfi = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put)
	begin
	  TASK_testplusargs___d446 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put)
	begin
	  TASK_testplusargs___d447 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put)
	begin
	  TASK_testplusargs___d448 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put)
	begin
	  v__h8601 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put &&
	  (TASK_testplusargs___d446 ||
	   TASK_testplusargs___d447 && TASK_testplusargs___d448))
	$write("[%10d", v__h8601, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put &&
	  (TASK_testplusargs___d446 ||
	   TASK_testplusargs___d447 && TASK_testplusargs___d448))
	$write("STAGE1: Writing RF[%d]:%h",
	       commit_rd_put[68:64],
	       commit_rd_put[63:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_commit_rd_put &&
	  (TASK_testplusargs___d446 ||
	   TASK_testplusargs___d447 && TASK_testplusargs___d448))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush)
	begin
	  TASK_testplusargs___d459 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush)
	begin
	  TASK_testplusargs___d460 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush)
	begin
	  TASK_testplusargs___d461 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush)
	begin
	  v__h8998 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush &&
	  (TASK_testplusargs___d459 ||
	   TASK_testplusargs___d460 && TASK_testplusargs___d461))
	$write("[%10d", v__h8998, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush &&
	  (TASK_testplusargs___d459 ||
	   TASK_testplusargs___d460 && TASK_testplusargs___d461))
	$write("STAGE1 : Received Flush. PC: %h ", ma_flush_newpc);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_flush &&
	  (TASK_testplusargs___d459 ||
	   TASK_testplusargs___d460 && TASK_testplusargs___d461))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize)
	begin
	  TASK_testplusargs___d2 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize)
	begin
	  TASK_testplusargs___d3 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize)
	begin
	  TASK_testplusargs___d4 = $test$plusargs("l1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize)
	begin
	  v__h2955 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize &&
	  (TASK_testplusargs___d2 ||
	   TASK_testplusargs___d3 && TASK_testplusargs___d4))
	$write("[%10d", v__h2955, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize &&
	  (TASK_testplusargs___d2 ||
	   TASK_testplusargs___d3 && TASK_testplusargs___d4))
	$write("STAGE1: Initializing the RF. Index: %d", rg_index);
    if (RST_N != `BSV_RESET_VALUE)
      if (rg_initialize &&
	  (TASK_testplusargs___d2 ||
	   TASK_testplusargs___d3 && TASK_testplusargs___d4))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt)
	begin
	  TASK_testplusargs___d17 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt)
	begin
	  TASK_testplusargs___d18 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt)
	begin
	  TASK_testplusargs___d19 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt)
	begin
	  v__h3340 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt &&
	  (TASK_testplusargs___d17 ||
	   TASK_testplusargs___d18 && TASK_testplusargs___d19))
	$write("[%10d", v__h3340, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt &&
	  (TASK_testplusargs___d17 ||
	   TASK_testplusargs___d18 && TASK_testplusargs___d19))
	$write("STAGE1 : Waiting for Interrupt. wr_interrupt: %b",
	       ma_interrupt_i);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_wait_for_interrupt &&
	  (TASK_testplusargs___d17 ||
	   TASK_testplusargs___d18 && TASK_testplusargs___d19))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65)
	begin
	  TASK_testplusargs___d91 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65)
	begin
	  TASK_testplusargs___d92 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65)
	begin
	  TASK_testplusargs___d93 = $test$plusargs("l1");
	  #0;
	end
    NOT_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_mem_ETC___d96 =
	!rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	(TASK_testplusargs___d91 ||
	 TASK_testplusargs___d92 && TASK_testplusargs___d93);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  !rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65)
	begin
	  v__h3536 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_mem_ETC___d96)
	$write("[%10d", v__h3536, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_mem_ETC___d96)
	$write("STAGE1 : Dropping Instruction from Cache");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_mem_ETC___d96)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d108 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d109 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d110 = $test$plusargs("l1");
	  #0;
	end
    TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d114 =
	(TASK_testplusargs___d108 ||
	 TASK_testplusargs___d109 && TASK_testplusargs___d110) &&
	rg_action;
    TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d115 =
	(TASK_testplusargs___d108 ||
	 TASK_testplusargs___d109 && TASK_testplusargs___d110) &&
	!rg_action;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h4359 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("[%10d", v__h4359, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("STAGE1 : rg_action: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d114)
	$write("None");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_08_OR_TASK_testplusargs_09_A_ETC___d115)
	$write("CheckPrev");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write(" Prev: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("PrevMeta { ", "instruction: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("'h%h", rg_prev[17:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write(", ", "epoch: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("'h%h", rg_prev[1:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write(" rg_discard:%b", rg_discard_lower);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d108 ||
	   TASK_testplusargs___d109 && TASK_testplusargs___d110))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d116 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d117 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d118 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h4531 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d116 ||
	   TASK_testplusargs___d117 && TASK_testplusargs___d118))
	$write("[%10d", v__h4531, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d116 ||
	   TASK_testplusargs___d117 && TASK_testplusargs___d118))
	$write("STAGE1: Decompressed: %h", _theResult_____4__h4464);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d116 ||
	   TASK_testplusargs___d117 && TASK_testplusargs___d118))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d168 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d169 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d170 = $test$plusargs("l3");
	  #0;
	end
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] == 2'd0;
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] == 2'd1;
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] == 2'd2;
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] != 2'd0 &&
	v_trigger_data1_0_wget[21:20] != 2'd1 &&
	v_trigger_data1_0_wget[21:20] != 2'd2;
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] != 2'd0 &&
	v_trigger_data1_0_wget[21:20] != 2'd1;
    TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195 =
	(TASK_testplusargs___d168 ||
	 TASK_testplusargs___d169 && TASK_testplusargs___d170) &&
	v_trigger_data1_0_wget[21:20] != 2'd0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h5120 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d168 ||
	   TASK_testplusargs___d169 && TASK_testplusargs___d170))
	$write("[%10d", v__h5120, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d168 ||
	   TASK_testplusargs___d169 && TASK_testplusargs___d170))
	$write("STAGE1 : Trigger[%2d] Data1: ", $signed(32'd0));
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("tagged MCONTROL ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("tagged ITRIGGER ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("tagged ETRIGGER ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("tagged NONE ", "");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("ETrigger { ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("'h%h", v_trigger_data1_0_wget[8:3]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("'h%h", v_trigger_data1_0_wget[2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("'h%h", v_trigger_data1_0_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d182)
	$write("'h%h", v_trigger_data1_0_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d188)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("ITrigger { ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("'h%h", v_trigger_data1_0_wget[8:3]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("'h%h", v_trigger_data1_0_wget[2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("'h%h", v_trigger_data1_0_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d180)
	$write("'h%h", v_trigger_data1_0_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d194)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("MControl { ", "load: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[19]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "store: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "execute: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[17]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "matched: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "chain: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[10]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[9:6]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "size: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[5:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "select: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d178)
	$write("'h%h", v_trigger_data1_0_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_68_OR_TASK_testplusargs_69_A_ETC___d195)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d168 ||
	   TASK_testplusargs___d169 && TASK_testplusargs___d170))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d205 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d206 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d207 = $test$plusargs("l3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h5546 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d205 ||
	   TASK_testplusargs___d206 && TASK_testplusargs___d207))
	$write("[%10d", v__h5546, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d205 ||
	   TASK_testplusargs___d206 && TASK_testplusargs___d207))
	$write("STAGE1 : Trigger[%2d] Data2: ",
	       $signed(32'd0),
	       "'h%h",
	       ma_trigger_data2_t[63:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d205 ||
	   TASK_testplusargs___d206 && TASK_testplusargs___d207))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d212 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d213 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d214 = $test$plusargs("l3");
	  #0;
	end
    TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d219 =
	(TASK_testplusargs___d212 ||
	 TASK_testplusargs___d213 && TASK_testplusargs___d214) &&
	ma_trigger_enable_t[0];
    TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d221 =
	(TASK_testplusargs___d212 ||
	 TASK_testplusargs___d213 && TASK_testplusargs___d214) &&
	!ma_trigger_enable_t[0];
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h5785 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d212 ||
	   TASK_testplusargs___d213 && TASK_testplusargs___d214))
	$write("[%10d", v__h5785, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d212 ||
	   TASK_testplusargs___d213 && TASK_testplusargs___d214))
	$write("STAGE1 : Trigger[%2d] Enable: ", $signed(32'd0));
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d219)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_12_OR_TASK_testplusargs_13_A_ETC___d221)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d212 ||
	   TASK_testplusargs___d213 && TASK_testplusargs___d214))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d222 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d223 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d224 = $test$plusargs("l3");
	  #0;
	end
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] == 2'd0;
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] == 2'd1;
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] == 2'd2;
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] != 2'd0 &&
	v_trigger_data1_1_wget[21:20] != 2'd1 &&
	v_trigger_data1_1_wget[21:20] != 2'd2;
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] != 2'd0;
    TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248 =
	(TASK_testplusargs___d222 ||
	 TASK_testplusargs___d223 && TASK_testplusargs___d224) &&
	v_trigger_data1_1_wget[21:20] != 2'd0 &&
	v_trigger_data1_1_wget[21:20] != 2'd1;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h6064 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d222 ||
	   TASK_testplusargs___d223 && TASK_testplusargs___d224))
	$write("[%10d", v__h6064, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d222 ||
	   TASK_testplusargs___d223 && TASK_testplusargs___d224))
	$write("STAGE1 : Trigger[%2d] Data1: ", $signed(32'd1));
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("tagged MCONTROL ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("tagged ITRIGGER ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("tagged ETRIGGER ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("tagged NONE ", "");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("ETrigger { ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("'h%h", v_trigger_data1_1_wget[8:3]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("'h%h", v_trigger_data1_1_wget[2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("'h%h", v_trigger_data1_1_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d236)
	$write("'h%h", v_trigger_data1_1_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d242)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("ITrigger { ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("'h%h", v_trigger_data1_1_wget[8:3]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("'h%h", v_trigger_data1_1_wget[2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("'h%h", v_trigger_data1_1_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d234)
	$write("'h%h", v_trigger_data1_1_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d248)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("MControl { ", "load: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[19]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "store: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "execute: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[17]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "user: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "machine: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "matched: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "chain: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[10]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "action_: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[9:6]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "size: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[5:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "select: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write(", ", "dmode: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d232)
	$write("'h%h", v_trigger_data1_1_wget[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_22_OR_TASK_testplusargs_23_A_ETC___d249)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d222 ||
	   TASK_testplusargs___d223 && TASK_testplusargs___d224))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d259 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d260 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d261 = $test$plusargs("l3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h6412 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d259 ||
	   TASK_testplusargs___d260 && TASK_testplusargs___d261))
	$write("[%10d", v__h6412, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d259 ||
	   TASK_testplusargs___d260 && TASK_testplusargs___d261))
	$write("STAGE1 : Trigger[%2d] Data2: ",
	       $signed(32'd1),
	       "'h%h",
	       ma_trigger_data2_t[127:64]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d259 ||
	   TASK_testplusargs___d260 && TASK_testplusargs___d261))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d266 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d267 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  TASK_testplusargs___d268 = $test$plusargs("l3");
	  #0;
	end
    TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d273 =
	(TASK_testplusargs___d266 ||
	 TASK_testplusargs___d267 && TASK_testplusargs___d268) &&
	ma_trigger_enable_t[1];
    TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d275 =
	(TASK_testplusargs___d266 ||
	 TASK_testplusargs___d267 && TASK_testplusargs___d268) &&
	!ma_trigger_enable_t[1];
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction)
	begin
	  v__h6581 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d266 ||
	   TASK_testplusargs___d267 && TASK_testplusargs___d268))
	$write("[%10d", v__h6581, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d266 ||
	   TASK_testplusargs___d267 && TASK_testplusargs___d268))
	$write("STAGE1 : Trigger[%2d] Enable: ", $signed(32'd1));
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d273)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  TASK_testplusargs_66_OR_TASK_testplusargs_67_A_ETC___d275)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  (TASK_testplusargs___d266 ||
	   TASK_testplusargs___d267 && TASK_testplusargs___d268))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d388 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d389 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d390 = $test$plusargs("l0");
	  #0;
	end
    NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393 =
	NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277 &&
	(TASK_testplusargs___d388 ||
	 TASK_testplusargs___d389 && TASK_testplusargs___d390);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  v__h7686 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("[%10d", v__h7686, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("STAGE1 : ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("TraceDump { ", "pc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("'h%h", rg_pc);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write(", ", "instruction: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("'h%h", final_instruction__h4155, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d393)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d395 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d396 = $test$plusargs("mstage1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  TASK_testplusargs___d397 = $test$plusargs("l1");
	  #0;
	end
    NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d400 =
	NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277 &&
	(TASK_testplusargs___d395 ||
	 TASK_testplusargs___d396 && TASK_testplusargs___d397);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d277)
	begin
	  v__h7835 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d400)
	$write("[%10d", v__h7835, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d400)
	$write("STAGE1 : compressed: %b perform_decode: %b curr_epoch: %b",
	       rg_eEpoch_6_CONCAT_rg_wEpoch_7_8_EQ_ff_memory__ETC___d65 &&
	       IF_NOT_rg_action_4_8_AND_rg_prev_1_BITS_1_TO_0_ETC___d124,
	       1'd1,
	       curr_epoch__h2865);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_process_instruction &&
	  NOT_IF_chk_interrupt_52_BIT_1_53_OR_ff_memory__ETC___d400)
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkstage1

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:15 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// rx_stage1_operands_deq_ena     O     1
// rx_stage1_meta_deq_ena         O     1
// rx_stage1_control_deq_ena      O     1
// tx_stage3_common_enq_ena       O     1
// tx_stage3_common_enq_data      O    70
// tx_stage3_type_enq_ena         O     1
// tx_stage3_type_enq_data        O    83
// rx_stage1_dump_deq_ena         O     1
// tx_stage3_dump_enq_ena         O     1
// tx_stage3_dump_enq_data        O    96
// memory_request_get             O   139
// RDY_memory_request_get         O     1 reg
// RDY_operand_fwding_put         O     1 const
// RDY_ma_update_wEpoch           O     1 const
// RDY_ma_csr_misa_c              O     1 const
// mv_delayed_output              O    65
// RDY_mv_delayed_output          O     1 const
// mv_redirection_fst             O    64
// RDY_mv_redirection_fst         O     1 const
// mv_redirection_snd             O     1
// RDY_mv_redirection_snd         O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// rx_stage1_operands_notEmpty_b  I     1 unused
// rx_stage1_operands_first_deq_rdy_b  I     1
// rx_stage1_operands_first_x     I   128
// rx_stage1_meta_notEmpty_b      I     1 unused
// rx_stage1_meta_first_deq_rdy_b  I     1
// rx_stage1_meta_first_x         I    65
// rx_stage1_control_notEmpty_b   I     1 unused
// rx_stage1_control_first_deq_rdy_b  I     1
// rx_stage1_control_first_x      I    66
// tx_stage3_common_notFull_b     I     1 unused
// tx_stage3_common_enq_rdy_b     I     1
// tx_stage3_type_notFull_b       I     1 unused
// tx_stage3_type_enq_rdy_b       I     1
// rx_stage1_dump_notEmpty_b      I     1 unused
// rx_stage1_dump_first_deq_rdy_b  I     1
// rx_stage1_dump_first_x         I    96
// tx_stage3_dump_notFull_b       I     1 unused
// tx_stage3_dump_enq_rdy_b       I     1
// operand_fwding_put             I    70
// ma_csr_misa_c_c                I     1
// ma_trigger_data1_t             I    44
// ma_trigger_data2_t             I   128
// ma_trigger_enable_t            I     2
// EN_operand_fwding_put          I     1
// EN_ma_update_wEpoch            I     1
// EN_ma_csr_misa_c               I     1
// EN_memory_request_get          I     1
//
// Combinational paths from inputs to outputs:
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> rx_stage1_operands_deq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> rx_stage1_meta_deq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> rx_stage1_control_deq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_common_enq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_common_enq_data
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_type_enq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_operands_first_x,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    ma_csr_misa_c_c,
//    ma_trigger_data1_t,
//    ma_trigger_data2_t,
//    ma_trigger_enable_t,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_type_enq_data
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> rx_stage1_dump_deq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_dump_enq_ena
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    rx_stage1_dump_first_x,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> tx_stage3_dump_enq_data
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_operands_first_x,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    ma_csr_misa_c_c,
//    ma_trigger_data1_t,
//    ma_trigger_data2_t,
//    ma_trigger_enable_t,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> mv_redirection_fst
//   (rx_stage1_operands_first_deq_rdy_b,
//    rx_stage1_operands_first_x,
//    rx_stage1_meta_first_deq_rdy_b,
//    rx_stage1_meta_first_x,
//    rx_stage1_control_first_deq_rdy_b,
//    rx_stage1_control_first_x,
//    tx_stage3_common_enq_rdy_b,
//    tx_stage3_type_enq_rdy_b,
//    rx_stage1_dump_first_deq_rdy_b,
//    tx_stage3_dump_enq_rdy_b,
//    operand_fwding_put,
//    ma_csr_misa_c_c,
//    ma_trigger_data1_t,
//    ma_trigger_data2_t,
//    ma_trigger_enable_t,
//    EN_operand_fwding_put,
//    EN_ma_csr_misa_c,
//    EN_memory_request_get) -> mv_redirection_snd
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkstage2(CLK,
		RST_N,

		rx_stage1_operands_notEmpty_b,

		rx_stage1_operands_first_deq_rdy_b,

		rx_stage1_operands_first_x,

		rx_stage1_operands_deq_ena,

		rx_stage1_meta_notEmpty_b,

		rx_stage1_meta_first_deq_rdy_b,

		rx_stage1_meta_first_x,

		rx_stage1_meta_deq_ena,

		rx_stage1_control_notEmpty_b,

		rx_stage1_control_first_deq_rdy_b,

		rx_stage1_control_first_x,

		rx_stage1_control_deq_ena,

		tx_stage3_common_notFull_b,

		tx_stage3_common_enq_rdy_b,

		tx_stage3_common_enq_ena,

		tx_stage3_common_enq_data,

		tx_stage3_type_notFull_b,

		tx_stage3_type_enq_rdy_b,

		tx_stage3_type_enq_ena,

		tx_stage3_type_enq_data,

		rx_stage1_dump_notEmpty_b,

		rx_stage1_dump_first_deq_rdy_b,

		rx_stage1_dump_first_x,

		rx_stage1_dump_deq_ena,

		tx_stage3_dump_notFull_b,

		tx_stage3_dump_enq_rdy_b,

		tx_stage3_dump_enq_ena,

		tx_stage3_dump_enq_data,

		EN_memory_request_get,
		memory_request_get,
		RDY_memory_request_get,

		operand_fwding_put,
		EN_operand_fwding_put,
		RDY_operand_fwding_put,

		EN_ma_update_wEpoch,
		RDY_ma_update_wEpoch,

		ma_csr_misa_c_c,
		EN_ma_csr_misa_c,
		RDY_ma_csr_misa_c,

		mv_delayed_output,
		RDY_mv_delayed_output,

		ma_trigger_data1_t,

		ma_trigger_data2_t,

		ma_trigger_enable_t,

		mv_redirection_fst,
		RDY_mv_redirection_fst,

		mv_redirection_snd,
		RDY_mv_redirection_snd);
  input  CLK;
  input  RST_N;

  // action method rx_stage1_operands_notEmpty
  input  rx_stage1_operands_notEmpty_b;

  // action method rx_stage1_operands_first_deq_rdy
  input  rx_stage1_operands_first_deq_rdy_b;

  // action method rx_stage1_operands_first
  input  [127 : 0] rx_stage1_operands_first_x;

  // value method rx_stage1_operands_deq_ena
  output rx_stage1_operands_deq_ena;

  // action method rx_stage1_meta_notEmpty
  input  rx_stage1_meta_notEmpty_b;

  // action method rx_stage1_meta_first_deq_rdy
  input  rx_stage1_meta_first_deq_rdy_b;

  // action method rx_stage1_meta_first
  input  [64 : 0] rx_stage1_meta_first_x;

  // value method rx_stage1_meta_deq_ena
  output rx_stage1_meta_deq_ena;

  // action method rx_stage1_control_notEmpty
  input  rx_stage1_control_notEmpty_b;

  // action method rx_stage1_control_first_deq_rdy
  input  rx_stage1_control_first_deq_rdy_b;

  // action method rx_stage1_control_first
  input  [65 : 0] rx_stage1_control_first_x;

  // value method rx_stage1_control_deq_ena
  output rx_stage1_control_deq_ena;

  // action method tx_stage3_common_notFull
  input  tx_stage3_common_notFull_b;

  // action method tx_stage3_common_enq_rdy
  input  tx_stage3_common_enq_rdy_b;

  // value method tx_stage3_common_enq_ena
  output tx_stage3_common_enq_ena;

  // value method tx_stage3_common_enq_data
  output [69 : 0] tx_stage3_common_enq_data;

  // action method tx_stage3_type_notFull
  input  tx_stage3_type_notFull_b;

  // action method tx_stage3_type_enq_rdy
  input  tx_stage3_type_enq_rdy_b;

  // value method tx_stage3_type_enq_ena
  output tx_stage3_type_enq_ena;

  // value method tx_stage3_type_enq_data
  output [82 : 0] tx_stage3_type_enq_data;

  // action method rx_stage1_dump_notEmpty
  input  rx_stage1_dump_notEmpty_b;

  // action method rx_stage1_dump_first_deq_rdy
  input  rx_stage1_dump_first_deq_rdy_b;

  // action method rx_stage1_dump_first
  input  [95 : 0] rx_stage1_dump_first_x;

  // value method rx_stage1_dump_deq_ena
  output rx_stage1_dump_deq_ena;

  // action method tx_stage3_dump_notFull
  input  tx_stage3_dump_notFull_b;

  // action method tx_stage3_dump_enq_rdy
  input  tx_stage3_dump_enq_rdy_b;

  // value method tx_stage3_dump_enq_ena
  output tx_stage3_dump_enq_ena;

  // value method tx_stage3_dump_enq_data
  output [95 : 0] tx_stage3_dump_enq_data;

  // actionvalue method memory_request_get
  input  EN_memory_request_get;
  output [138 : 0] memory_request_get;
  output RDY_memory_request_get;

  // action method operand_fwding_put
  input  [69 : 0] operand_fwding_put;
  input  EN_operand_fwding_put;
  output RDY_operand_fwding_put;

  // action method ma_update_wEpoch
  input  EN_ma_update_wEpoch;
  output RDY_ma_update_wEpoch;

  // action method ma_csr_misa_c
  input  ma_csr_misa_c_c;
  input  EN_ma_csr_misa_c;
  output RDY_ma_csr_misa_c;

  // value method mv_delayed_output
  output [64 : 0] mv_delayed_output;
  output RDY_mv_delayed_output;

  // action method ma_trigger_data1
  input  [43 : 0] ma_trigger_data1_t;

  // action method ma_trigger_data2
  input  [127 : 0] ma_trigger_data2_t;

  // action method ma_trigger_enable
  input  [1 : 0] ma_trigger_enable_t;

  // value method mv_redirection_fst
  output [63 : 0] mv_redirection_fst;
  output RDY_mv_redirection_fst;

  // value method mv_redirection_snd
  output mv_redirection_snd;
  output RDY_mv_redirection_snd;

  // signals for module outputs
  wire [138 : 0] memory_request_get;
  wire [95 : 0] tx_stage3_dump_enq_data;
  wire [82 : 0] tx_stage3_type_enq_data;
  wire [69 : 0] tx_stage3_common_enq_data;
  wire [64 : 0] mv_delayed_output;
  wire [63 : 0] mv_redirection_fst;
  wire RDY_ma_csr_misa_c,
       RDY_ma_update_wEpoch,
       RDY_memory_request_get,
       RDY_mv_delayed_output,
       RDY_mv_redirection_fst,
       RDY_mv_redirection_snd,
       RDY_operand_fwding_put,
       mv_redirection_snd,
       rx_stage1_control_deq_ena,
       rx_stage1_dump_deq_ena,
       rx_stage1_meta_deq_ena,
       rx_stage1_operands_deq_ena,
       tx_stage3_common_enq_ena,
       tx_stage3_dump_enq_ena,
       tx_stage3_type_enq_ena;

  // inlined wires
  reg [21 : 0] v_trigger_data1_0_wget, v_trigger_data1_1_wget;
  wire [82 : 0] ff_stage3_type_w_data_wget;
  wire [69 : 0] ff_stage3_common_w_data_wget;
  wire [64 : 0] ff_stage1_meta_w_data_wget, wr_redirection_wget;
  wire ff_stage1_operands_w_ena_whas, ff_stage3_common_w_ena_whas;

  // register rg_eEpoch
  reg rg_eEpoch;
  wire rg_eEpoch_D_IN, rg_eEpoch_EN;

  // register rg_loadreserved_addr
  reg [32 : 0] rg_loadreserved_addr;
  wire [32 : 0] rg_loadreserved_addr_D_IN;
  wire rg_loadreserved_addr_EN;

  // register rg_wEpoch
  reg rg_wEpoch;
  wire rg_wEpoch_D_IN, rg_wEpoch_EN;

  // ports of submodule alu
  reg [63 : 0] alu_inputs_op3;
  reg [1 : 0] alu_inputs_memaccess;
  wire [137 : 0] alu_inputs;
  wire [127 : 0] alu_inputs_tdata2;
  wire [64 : 0] alu_mv_delayed_output;
  wire [63 : 0] alu_inputs_imm_value, alu_inputs_op1, alu_inputs_op2;
  wire [43 : 0] alu_inputs_tdata1;
  wire [3 : 0] alu_inputs_fn, alu_inputs_inst_type;
  wire [2 : 0] alu_inputs_funct3;
  wire [1 : 0] alu_inputs_lpc, alu_inputs_tenable;
  wire alu_EN_inputs, alu_inputs_misa_c, alu_inputs_word32;

  // ports of submodule ff_memory_request
  wire [138 : 0] ff_memory_request_D_IN, ff_memory_request_D_OUT;
  wire ff_memory_request_CLR,
       ff_memory_request_DEQ,
       ff_memory_request_EMPTY_N,
       ff_memory_request_ENQ,
       ff_memory_request_FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_fetch_execute_pass,
       CAN_FIRE_ma_csr_misa_c,
       CAN_FIRE_ma_trigger_data1,
       CAN_FIRE_ma_trigger_data2,
       CAN_FIRE_ma_trigger_enable,
       CAN_FIRE_ma_update_wEpoch,
       CAN_FIRE_memory_request_get,
       CAN_FIRE_operand_fwding_put,
       CAN_FIRE_rx_stage1_control_first,
       CAN_FIRE_rx_stage1_control_first_deq_rdy,
       CAN_FIRE_rx_stage1_control_notEmpty,
       CAN_FIRE_rx_stage1_dump_first,
       CAN_FIRE_rx_stage1_dump_first_deq_rdy,
       CAN_FIRE_rx_stage1_dump_notEmpty,
       CAN_FIRE_rx_stage1_meta_first,
       CAN_FIRE_rx_stage1_meta_first_deq_rdy,
       CAN_FIRE_rx_stage1_meta_notEmpty,
       CAN_FIRE_rx_stage1_operands_first,
       CAN_FIRE_rx_stage1_operands_first_deq_rdy,
       CAN_FIRE_rx_stage1_operands_notEmpty,
       CAN_FIRE_tx_stage3_common_enq_rdy,
       CAN_FIRE_tx_stage3_common_notFull,
       CAN_FIRE_tx_stage3_dump_enq_rdy,
       CAN_FIRE_tx_stage3_dump_notFull,
       CAN_FIRE_tx_stage3_type_enq_rdy,
       CAN_FIRE_tx_stage3_type_notFull,
       WILL_FIRE_RL_fetch_execute_pass,
       WILL_FIRE_ma_csr_misa_c,
       WILL_FIRE_ma_trigger_data1,
       WILL_FIRE_ma_trigger_data2,
       WILL_FIRE_ma_trigger_enable,
       WILL_FIRE_ma_update_wEpoch,
       WILL_FIRE_memory_request_get,
       WILL_FIRE_operand_fwding_put,
       WILL_FIRE_rx_stage1_control_first,
       WILL_FIRE_rx_stage1_control_first_deq_rdy,
       WILL_FIRE_rx_stage1_control_notEmpty,
       WILL_FIRE_rx_stage1_dump_first,
       WILL_FIRE_rx_stage1_dump_first_deq_rdy,
       WILL_FIRE_rx_stage1_dump_notEmpty,
       WILL_FIRE_rx_stage1_meta_first,
       WILL_FIRE_rx_stage1_meta_first_deq_rdy,
       WILL_FIRE_rx_stage1_meta_notEmpty,
       WILL_FIRE_rx_stage1_operands_first,
       WILL_FIRE_rx_stage1_operands_first_deq_rdy,
       WILL_FIRE_rx_stage1_operands_notEmpty,
       WILL_FIRE_tx_stage3_common_enq_rdy,
       WILL_FIRE_tx_stage3_common_notFull,
       WILL_FIRE_tx_stage3_dump_enq_rdy,
       WILL_FIRE_tx_stage3_dump_notFull,
       WILL_FIRE_tx_stage3_type_enq_rdy,
       WILL_FIRE_tx_stage3_type_notFull;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d30;
  reg TASK_testplusargs___d31;
  reg TASK_testplusargs___d32;
  reg [63 : 0] v__h3163;
  reg TASK_testplusargs___d42;
  reg TASK_testplusargs___d43;
  reg TASK_testplusargs___d44;
  reg [63 : 0] v__h3348;
  reg TASK_testplusargs___d54;
  reg TASK_testplusargs___d55;
  reg TASK_testplusargs___d56;
  reg [63 : 0] v__h3537;
  reg TASK_testplusargs___d126;
  reg TASK_testplusargs___d127;
  reg TASK_testplusargs___d128;
  reg [63 : 0] v__h3898;
  reg TASK_testplusargs___d138;
  reg TASK_testplusargs___d139;
  reg TASK_testplusargs___d140;
  reg [63 : 0] v__h4078;
  reg TASK_testplusargs___d164;
  reg TASK_testplusargs___d165;
  reg TASK_testplusargs___d166;
  reg [63 : 0] v__h4298;
  reg TASK_testplusargs___d176;
  reg TASK_testplusargs___d177;
  reg TASK_testplusargs___d178;
  reg [63 : 0] v__h4485;
  reg TASK_testplusargs___d239;
  reg TASK_testplusargs___d240;
  reg TASK_testplusargs___d241;
  reg [63 : 0] v__h6283;
  reg TASK_testplusargs___d294;
  reg TASK_testplusargs___d295;
  reg TASK_testplusargs___d296;
  reg [63 : 0] v__h6977;
  reg TASK_testplusargs___d311;
  reg TASK_testplusargs___d312;
  reg TASK_testplusargs___d313;
  reg [63 : 0] v__h7230;
  reg TASK_testplusargs___d391;
  reg TASK_testplusargs___d392;
  reg TASK_testplusargs___d393;
  reg [63 : 0] v__h6617;
  reg TASK_testplusargs___d470;
  reg TASK_testplusargs___d471;
  reg TASK_testplusargs___d472;
  reg [63 : 0] v__h9106;
  reg IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d299;
  reg IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d316;
  reg TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d323;
  reg TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d330;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d65;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d67;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d69;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d71;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d73;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d75;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d77;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d79;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d95;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d105;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d107;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d109;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d115;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d123;
  reg TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d125;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d147;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d149;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d153;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d155;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d157;
  reg TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d163;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d247;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d249;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d252;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d254;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d256;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d262;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d267;
  reg TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d269;
  reg IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d302;
  reg IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d319;
  reg NOT_IF_ff_stage1_control_w_data_whas__70_THEN__ETC___d396;
  // synopsys translate_on

  // remaining internal signals
  reg [82 : 0] IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d388;
  reg [63 : 0] _op2__h3087;
  reg [21 : 0] CASE_v_trigger_data1_0wget_BITS_21_TO_20_0_v__ETC__q8,
	       CASE_v_trigger_data1_1wget_BITS_21_TO_20_0_v__ETC__q7;
  reg [1 : 0] CASE_IF_ff_stage3_type_w_data_whas__23_THEN_IF_ETC__q6,
	      CASE_ff_memory_requestD_OUT_BITS_10_TO_9_0_ff_ETC__q2,
	      CASE_rx_stage1_meta_first_x_BITS_42_TO_41_0_rx_ETC__q1,
	      IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356,
	      IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103,
	      IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435;
  wire [63 : 0] SEXT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff__ETC___d203,
		_theResult_____1_snd_aluresult__h7454,
		op1__h3084,
		op2__h3085,
		rd__h4543,
		rx_stage1_control_first_x_BITS_63_TO_0__q5,
		s3regular_rdvalue__h7827,
		s3system_rs1_imm__h7842,
		x1_avValue_snd_aluresult__h7460;
  wire [31 : 0] ff_stage1_meta_w_datawget_BITS_40_TO_9__q4;
  wire [6 : 0] ff_stage1_meta_w_datawget_BITS_8_TO_2__q3;
  wire [4 : 0] rdaddr__h4542, x__h6827;
  wire [1 : 0] IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305,
	       IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d340,
	       IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341,
	       IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346,
	       IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d339,
	       IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d344,
	       curr_epoch__h1856;
  wire IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273,
       IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d186,
       IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d188,
       NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195,
       NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292,
       NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309,
       NOT_alu_inputs_45_BITS_38_TO_7_88_EQ_rg_loadre_ETC___d336,
       v_trigger_enable_0_whas_AND_ff_stage1_dump_w_r_ETC___d21;

  // action method rx_stage1_operands_notEmpty
  assign CAN_FIRE_rx_stage1_operands_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage1_operands_notEmpty = 1'd1 ;

  // action method rx_stage1_operands_first_deq_rdy
  assign CAN_FIRE_rx_stage1_operands_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage1_operands_first_deq_rdy = 1'd1 ;

  // action method rx_stage1_operands_first
  assign CAN_FIRE_rx_stage1_operands_first = 1'd1 ;
  assign WILL_FIRE_rx_stage1_operands_first = 1'd1 ;

  // value method rx_stage1_operands_deq_ena
  assign rx_stage1_operands_deq_ena = ff_stage1_operands_w_ena_whas ;

  // action method rx_stage1_meta_notEmpty
  assign CAN_FIRE_rx_stage1_meta_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage1_meta_notEmpty = 1'd1 ;

  // action method rx_stage1_meta_first_deq_rdy
  assign CAN_FIRE_rx_stage1_meta_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage1_meta_first_deq_rdy = 1'd1 ;

  // action method rx_stage1_meta_first
  assign CAN_FIRE_rx_stage1_meta_first = 1'd1 ;
  assign WILL_FIRE_rx_stage1_meta_first = 1'd1 ;

  // value method rx_stage1_meta_deq_ena
  assign rx_stage1_meta_deq_ena = ff_stage1_operands_w_ena_whas ;

  // action method rx_stage1_control_notEmpty
  assign CAN_FIRE_rx_stage1_control_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage1_control_notEmpty = 1'd1 ;

  // action method rx_stage1_control_first_deq_rdy
  assign CAN_FIRE_rx_stage1_control_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage1_control_first_deq_rdy = 1'd1 ;

  // action method rx_stage1_control_first
  assign CAN_FIRE_rx_stage1_control_first = 1'd1 ;
  assign WILL_FIRE_rx_stage1_control_first = 1'd1 ;

  // value method rx_stage1_control_deq_ena
  assign rx_stage1_control_deq_ena = ff_stage1_operands_w_ena_whas ;

  // action method tx_stage3_common_notFull
  assign CAN_FIRE_tx_stage3_common_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage3_common_notFull = 1'd1 ;

  // action method tx_stage3_common_enq_rdy
  assign CAN_FIRE_tx_stage3_common_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage3_common_enq_rdy = 1'd1 ;

  // value method tx_stage3_common_enq_ena
  assign tx_stage3_common_enq_ena = ff_stage3_common_w_ena_whas ;

  // value method tx_stage3_common_enq_data
  assign tx_stage3_common_enq_data = ff_stage3_common_w_data_wget ;

  // action method tx_stage3_type_notFull
  assign CAN_FIRE_tx_stage3_type_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage3_type_notFull = 1'd1 ;

  // action method tx_stage3_type_enq_rdy
  assign CAN_FIRE_tx_stage3_type_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage3_type_enq_rdy = 1'd1 ;

  // value method tx_stage3_type_enq_ena
  assign tx_stage3_type_enq_ena = ff_stage3_common_w_ena_whas ;

  // value method tx_stage3_type_enq_data
  assign tx_stage3_type_enq_data =
	     (ff_stage3_common_w_ena_whas &&
	      ff_stage3_type_w_data_wget[82:81] == 2'd0) ?
	       { 2'd0,
		 13'b0101010101010 /* unspecified value */ ,
		 CASE_IF_ff_stage3_type_w_data_whas__23_THEN_IF_ETC__q6,
		 ff_stage3_type_w_data_wget[65:0] } :
	       { (ff_stage3_common_w_ena_whas &&
		  ff_stage3_type_w_data_wget[82:81] == 2'd1) ?
		   2'd1 :
		   ((ff_stage3_common_w_ena_whas &&
		     ff_stage3_type_w_data_wget[82:81] == 2'd2) ?
		      2'd2 :
		      2'd3),
		 ff_stage3_type_w_data_wget[80:0] } ;

  // action method rx_stage1_dump_notEmpty
  assign CAN_FIRE_rx_stage1_dump_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage1_dump_notEmpty = 1'd1 ;

  // action method rx_stage1_dump_first_deq_rdy
  assign CAN_FIRE_rx_stage1_dump_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage1_dump_first_deq_rdy = 1'd1 ;

  // action method rx_stage1_dump_first
  assign CAN_FIRE_rx_stage1_dump_first = 1'd1 ;
  assign WILL_FIRE_rx_stage1_dump_first = 1'd1 ;

  // value method rx_stage1_dump_deq_ena
  assign rx_stage1_dump_deq_ena = ff_stage1_operands_w_ena_whas ;

  // action method tx_stage3_dump_notFull
  assign CAN_FIRE_tx_stage3_dump_notFull = 1'd1 ;
  assign WILL_FIRE_tx_stage3_dump_notFull = 1'd1 ;

  // action method tx_stage3_dump_enq_rdy
  assign CAN_FIRE_tx_stage3_dump_enq_rdy = 1'd1 ;
  assign WILL_FIRE_tx_stage3_dump_enq_rdy = 1'd1 ;

  // value method tx_stage3_dump_enq_ena
  assign tx_stage3_dump_enq_ena = ff_stage3_common_w_ena_whas ;

  // value method tx_stage3_dump_enq_data
  assign tx_stage3_dump_enq_data = rx_stage1_dump_first_x ;

  // actionvalue method memory_request_get
  assign memory_request_get =
	     { ff_memory_request_D_OUT[138:11],
	       CASE_ff_memory_requestD_OUT_BITS_10_TO_9_0_ff_ETC__q2,
	       ff_memory_request_D_OUT[8:0] } ;
  assign RDY_memory_request_get = ff_memory_request_EMPTY_N ;
  assign CAN_FIRE_memory_request_get = ff_memory_request_EMPTY_N ;
  assign WILL_FIRE_memory_request_get = EN_memory_request_get ;

  // action method operand_fwding_put
  assign RDY_operand_fwding_put = 1'd1 ;
  assign CAN_FIRE_operand_fwding_put = 1'd1 ;
  assign WILL_FIRE_operand_fwding_put = EN_operand_fwding_put ;

  // action method ma_update_wEpoch
  assign RDY_ma_update_wEpoch = 1'd1 ;
  assign CAN_FIRE_ma_update_wEpoch = 1'd1 ;
  assign WILL_FIRE_ma_update_wEpoch = EN_ma_update_wEpoch ;

  // action method ma_csr_misa_c
  assign RDY_ma_csr_misa_c = 1'd1 ;
  assign CAN_FIRE_ma_csr_misa_c = 1'd1 ;
  assign WILL_FIRE_ma_csr_misa_c = EN_ma_csr_misa_c ;

  // value method mv_delayed_output
  assign mv_delayed_output = alu_mv_delayed_output ;
  assign RDY_mv_delayed_output = 1'd1 ;

  // action method ma_trigger_data1
  assign CAN_FIRE_ma_trigger_data1 = 1'd1 ;
  assign WILL_FIRE_ma_trigger_data1 = 1'd1 ;

  // action method ma_trigger_data2
  assign CAN_FIRE_ma_trigger_data2 = 1'd1 ;
  assign WILL_FIRE_ma_trigger_data2 = 1'd1 ;

  // action method ma_trigger_enable
  assign CAN_FIRE_ma_trigger_enable = 1'd1 ;
  assign WILL_FIRE_ma_trigger_enable = 1'd1 ;

  // value method mv_redirection_fst
  assign mv_redirection_fst = wr_redirection_wget[64:1] ;
  assign RDY_mv_redirection_fst = 1'd1 ;

  // value method mv_redirection_snd
  assign mv_redirection_snd =
	     ff_stage3_common_w_ena_whas && wr_redirection_wget[0] ;
  assign RDY_mv_redirection_snd = 1'd1 ;

  // submodule alu
  mkalu alu(.CLK(CLK),
	    .RST_N(RST_N),
	    .inputs_fn(alu_inputs_fn),
	    .inputs_funct3(alu_inputs_funct3),
	    .inputs_imm_value(alu_inputs_imm_value),
	    .inputs_inst_type(alu_inputs_inst_type),
	    .inputs_lpc(alu_inputs_lpc),
	    .inputs_memaccess(alu_inputs_memaccess),
	    .inputs_misa_c(alu_inputs_misa_c),
	    .inputs_op1(alu_inputs_op1),
	    .inputs_op2(alu_inputs_op2),
	    .inputs_op3(alu_inputs_op3),
	    .inputs_tdata1(alu_inputs_tdata1),
	    .inputs_tdata2(alu_inputs_tdata2),
	    .inputs_tenable(alu_inputs_tenable),
	    .inputs_word32(alu_inputs_word32),
	    .EN_inputs(alu_EN_inputs),
	    .inputs(alu_inputs),
	    .RDY_inputs(),
	    .mv_delayed_output(alu_mv_delayed_output),
	    .RDY_mv_delayed_output());

  // submodule ff_memory_request
  FIFOL1 #(.width(32'd139)) ff_memory_request(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(ff_memory_request_D_IN),
					      .ENQ(ff_memory_request_ENQ),
					      .DEQ(ff_memory_request_DEQ),
					      .CLR(ff_memory_request_CLR),
					      .D_OUT(ff_memory_request_D_OUT),
					      .FULL_N(ff_memory_request_FULL_N),
					      .EMPTY_N(ff_memory_request_EMPTY_N));

  // rule RL_fetch_execute_pass
  assign CAN_FIRE_RL_fetch_execute_pass =
	     rx_stage1_meta_first_deq_rdy_b &&
	     rx_stage1_control_first_deq_rdy_b &&
	     EN_ma_csr_misa_c &&
	     v_trigger_enable_0_whas_AND_ff_stage1_dump_w_r_ETC___d21 ;
  assign WILL_FIRE_RL_fetch_execute_pass = CAN_FIRE_RL_fetch_execute_pass ;

  // inlined wires
  assign ff_stage1_operands_w_ena_whas =
	     WILL_FIRE_RL_fetch_execute_pass &&
	     (NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 ||
	      !IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273) ;
  assign ff_stage1_meta_w_data_wget =
	     { rx_stage1_meta_first_x[64:43],
	       CASE_rx_stage1_meta_first_x_BITS_42_TO_41_0_rx_ETC__q1,
	       rx_stage1_meta_first_x[40:0] } ;
  assign ff_stage3_common_w_ena_whas =
	     WILL_FIRE_RL_fetch_execute_pass &&
	     IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 ;
  assign ff_stage3_common_w_data_wget =
	     { rx_stage1_control_first_x[63:0],
	       ff_stage1_meta_w_data_wget[54:50],
	       rg_wEpoch } ;
  assign ff_stage3_type_w_data_wget =
	     (IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 !=
	      2'd2 &&
	      IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 !=
	      2'd1 &&
	      IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 !=
	      2'd3) ?
	       { 2'd0,
		 13'b0101010101010 /* unspecified value */ ,
		 IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356,
		 alu_inputs[70:7],
		 ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[1:0] } :
	       IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d388 ;
  assign wr_redirection_wget = { alu_inputs[70:7], alu_inputs[0] } ;
  always@(ma_trigger_data1_t)
  begin
    case (ma_trigger_data1_t[21:20])
      2'd0, 2'd1, 2'd2: v_trigger_data1_0_wget = ma_trigger_data1_t[21:0];
      2'd3:
	  v_trigger_data1_0_wget =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(ma_trigger_data1_t)
  begin
    case (ma_trigger_data1_t[43:42])
      2'd0, 2'd1, 2'd2: v_trigger_data1_1_wget = ma_trigger_data1_t[43:22];
      2'd3:
	  v_trigger_data1_1_wget =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end

  // register rg_eEpoch
  assign rg_eEpoch_D_IN = ~rg_eEpoch ;
  assign rg_eEpoch_EN =
	     WILL_FIRE_RL_fetch_execute_pass &&
	     IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	     alu_inputs[0] ;

  // register rg_loadreserved_addr
  assign rg_loadreserved_addr_D_IN =
	     { x__h6827 == 5'b00101 &&
	       IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 ==
	       2'd3,
	       alu_inputs[38:7] } ;
  assign rg_loadreserved_addr_EN =
	     WILL_FIRE_RL_fetch_execute_pass &&
	     IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	     ff_stage1_meta_w_data_wget[46:43] == 4'd1 ;

  // register rg_wEpoch
  assign rg_wEpoch_D_IN = ~rg_wEpoch ;
  assign rg_wEpoch_EN = EN_ma_update_wEpoch ;

  // submodule alu
  assign alu_inputs_fn = ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[6:3] ;
  assign alu_inputs_funct3 = ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[2:0] ;
  assign alu_inputs_imm_value =
	     SEXT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff__ETC___d203 ;
  assign alu_inputs_inst_type = ff_stage1_meta_w_data_wget[46:43] ;
  assign alu_inputs_lpc = rx_stage1_control_first_x_BITS_63_TO_0__q5[1:0] ;
  always@(IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103)
  begin
    case (IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103)
      2'd0, 2'd1:
	  alu_inputs_memaccess =
	      IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103;
      2'd2: alu_inputs_memaccess = 2'd3;
      2'd3: alu_inputs_memaccess = 2'd2;
    endcase
  end
  assign alu_inputs_misa_c = ma_csr_misa_c_c ;
  assign alu_inputs_op1 =
	     ff_stage1_meta_w_data_wget[49] ?
	       rx_stage1_control_first_x[63:0] :
	       op1__h3084 ;
  assign alu_inputs_op2 = _op2__h3087 ;
  always@(ff_stage1_meta_w_data_wget or
	  rx_stage1_control_first_x or op1__h3084)
  begin
    case (ff_stage1_meta_w_data_wget[46:43])
      4'd1, 4'd4: alu_inputs_op3 = op1__h3084;
      default: alu_inputs_op3 = rx_stage1_control_first_x[63:0];
    endcase
  end
  assign alu_inputs_tdata1 =
	     { CASE_v_trigger_data1_1wget_BITS_21_TO_20_0_v__ETC__q7,
	       CASE_v_trigger_data1_0wget_BITS_21_TO_20_0_v__ETC__q8 } ;
  assign alu_inputs_tdata2 = ma_trigger_data2_t ;
  assign alu_inputs_tenable = ma_trigger_enable_t ;
  assign alu_inputs_word32 = ff_stage1_meta_w_data_wget[1] ;
  assign alu_EN_inputs = CAN_FIRE_RL_fetch_execute_pass ;

  // submodule ff_memory_request
  assign ff_memory_request_D_IN =
	     { alu_inputs[70:7],
	       _op2__h3087,
	       IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356,
	       ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[2:0],
	       rg_wEpoch,
	       x__h6827 } ;
  assign ff_memory_request_ENQ =
	     WILL_FIRE_RL_fetch_execute_pass &&
	     IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	     IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 ==
	     2'd0 &&
	     IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346 !=
	     2'd2 ;
  assign ff_memory_request_DEQ = EN_memory_request_get ;
  assign ff_memory_request_CLR = EN_ma_update_wEpoch ;

  // remaining internal signals
  assign IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 =
	     (x__h6827 == 5'b00101 &&
	      IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 ==
	      2'd3) ?
	       2'd0 :
	       IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 ;
  assign IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d340 =
	     (x__h6827 == 5'b00111 &&
	      IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 ==
	      2'd3) ?
	       IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d339 :
	       alu_inputs[136:135] ;
  assign IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 =
	     (ff_stage1_meta_w_data_wget[46:43] == 4'd1) ?
	       IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d340 :
	       alu_inputs[136:135] ;
  assign IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346 =
	     (ff_stage1_meta_w_data_wget[46:43] == 4'd1) ?
	       ((x__h6827 == 5'b00111 &&
		 IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 ==
		 2'd3) ?
		  IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d344 :
		  IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305) :
	       IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 ;
  assign IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 =
	     rx_stage1_control_first_x[65:64] == curr_epoch__h1856 ;
  assign IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d186 =
	     ff_stage1_meta_w_data_wget[64:60] == rdaddr__h4542 ;
  assign IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d188 =
	     ff_stage1_meta_w_data_wget[59:55] == rdaddr__h4542 ;
  assign IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d339 =
	     (rg_loadreserved_addr[32] &&
	      NOT_alu_inputs_45_BITS_38_TO_7_88_EQ_rg_loadre_ETC___d336) ?
	       2'd2 :
	       (rg_loadreserved_addr[32] ? alu_inputs[136:135] : 2'd2) ;
  assign IF_rg_loadreserved_addr_21_BIT_32_22_AND_NOT_a_ETC___d344 =
	     (rg_loadreserved_addr[32] &&
	      NOT_alu_inputs_45_BITS_38_TO_7_88_EQ_rg_loadre_ETC___d336) ?
	       IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 :
	       (rg_loadreserved_addr[32] ?
		  2'd1 :
		  IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305) ;
  assign NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 =
	     !IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d186 &&
	     !IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d188 ||
	     EN_operand_fwding_put && operand_fwding_put[0] ||
	     rdaddr__h4542 == 5'd0 ;
  assign NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292 =
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	     ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	     x__h6827 == 5'b00101 &&
	     IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 ==
	     2'd3 ;
  assign NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309 =
	     NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	     ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	     x__h6827 == 5'b00111 &&
	     IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 ==
	     2'd3 ;
  assign NOT_alu_inputs_45_BITS_38_TO_7_88_EQ_rg_loadre_ETC___d336 =
	     alu_inputs[38:7] != rg_loadreserved_addr[31:0] ;
  assign SEXT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff__ETC___d203 =
	     { {32{ff_stage1_meta_w_datawget_BITS_40_TO_9__q4[31]}},
	       ff_stage1_meta_w_datawget_BITS_40_TO_9__q4 } ;
  assign _theResult_____1_snd_aluresult__h7454 =
	     (NOT_alu_inputs_45_BITS_38_TO_7_88_EQ_rg_loadre_ETC___d336 ||
	      !rg_loadreserved_addr[32]) ?
	       64'd1 :
	       alu_inputs[134:71] ;
  assign curr_epoch__h1856 = { rg_eEpoch, rg_wEpoch } ;
  assign ff_stage1_meta_w_datawget_BITS_40_TO_9__q4 =
	     ff_stage1_meta_w_data_wget[40:9] ;
  assign ff_stage1_meta_w_datawget_BITS_8_TO_2__q3 =
	     ff_stage1_meta_w_data_wget[8:2] ;
  assign op1__h3084 =
	     IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d186 ?
	       rd__h4543 :
	       rx_stage1_operands_first_x[127:64] ;
  assign op2__h3085 =
	     IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d188 ?
	       rd__h4543 :
	       rx_stage1_operands_first_x[63:0] ;
  assign rd__h4543 =
	     EN_operand_fwding_put ? operand_fwding_put[64:1] : 64'd0 ;
  assign rdaddr__h4542 =
	     EN_operand_fwding_put ? operand_fwding_put[69:65] : 5'd0 ;
  assign rx_stage1_control_first_x_BITS_63_TO_0__q5 =
	     rx_stage1_control_first_x[63:0] ;
  assign s3regular_rdvalue__h7827 =
	     (ff_stage1_meta_w_data_wget[46:43] == 4'd1) ?
	       x1_avValue_snd_aluresult__h7460 :
	       alu_inputs[134:71] ;
  assign s3system_rs1_imm__h7842 =
	     ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[2] ?
	       { 59'd0, ff_stage1_meta_w_datawget_BITS_40_TO_9__q4[16:12] } :
	       s3regular_rdvalue__h7827 ;
  assign v_trigger_enable_0_whas_AND_ff_stage1_dump_w_r_ETC___d21 =
	     rx_stage1_dump_first_deq_rdy_b &&
	     rx_stage1_operands_first_deq_rdy_b &&
	     tx_stage3_common_enq_rdy_b &&
	     tx_stage3_type_enq_rdy_b &&
	     tx_stage3_dump_enq_rdy_b &&
	     ff_memory_request_FULL_N ;
  assign x1_avValue_snd_aluresult__h7460 =
	     (x__h6827 == 5'b00111 &&
	      IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 ==
	      2'd3) ?
	       _theResult_____1_snd_aluresult__h7454 :
	       alu_inputs[134:71] ;
  assign x__h6827 =
	     { ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[0],
	       ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[6:3] } ;
  always@(rx_stage1_meta_first_x)
  begin
    case (rx_stage1_meta_first_x[42:41])
      2'd0, 2'd1, 2'd3:
	  CASE_rx_stage1_meta_first_x_BITS_42_TO_41_0_rx_ETC__q1 =
	      rx_stage1_meta_first_x[42:41];
      2'd2: CASE_rx_stage1_meta_first_x_BITS_42_TO_41_0_rx_ETC__q1 = 2'd2;
    endcase
  end
  always@(ff_memory_request_D_OUT)
  begin
    case (ff_memory_request_D_OUT[10:9])
      2'd0, 2'd1, 2'd3:
	  CASE_ff_memory_requestD_OUT_BITS_10_TO_9_0_ff_ETC__q2 =
	      ff_memory_request_D_OUT[10:9];
      2'd2: CASE_ff_memory_requestD_OUT_BITS_10_TO_9_0_ff_ETC__q2 = 2'd2;
    endcase
  end
  always@(ff_stage1_meta_w_data_wget)
  begin
    case (ff_stage1_meta_w_data_wget[42:41])
      2'd0, 2'd1:
	  IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 =
	      ff_stage1_meta_w_data_wget[42:41];
      2'd2: IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 = 2'd3;
      2'd3: IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 = 2'd2;
    endcase
  end
  always@(IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346)
  begin
    case (IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346)
      2'd0, 2'd1:
	  IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356 =
	      IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d346;
      2'd2: IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356 = 2'd3;
      2'd3: IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d356 = 2'd2;
    endcase
  end
  always@(ff_stage1_meta_w_data_wget or
	  op2__h3085 or
	  SEXT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff__ETC___d203)
  begin
    case (ff_stage1_meta_w_data_wget[48:47])
      2'd0: _op2__h3087 = op2__h3085;
      2'd1:
	  _op2__h3087 =
	      SEXT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff__ETC___d203;
      2'd2: _op2__h3087 = 64'd4;
      2'd3: _op2__h3087 = 64'd2;
    endcase
  end
  always@(IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341 or
	  s3system_rs1_imm__h7842 or
	  rx_stage1_control_first_x_BITS_63_TO_0__q5 or
	  ff_stage1_meta_w_datawget_BITS_40_TO_9__q4 or
	  ff_stage1_meta_w_datawget_BITS_8_TO_2__q3 or
	  s3regular_rdvalue__h7827 or alu_inputs)
  begin
    case (IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341)
      2'd2:
	  IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d388 =
	      { IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d341,
		16'b1010101010101010 /* unspecified value */ ,
		s3regular_rdvalue__h7827,
		!alu_inputs[137] };
      2'd3:
	  IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d388 =
	      { 2'd1,
		11'b01010101010 /* unspecified value */ ,
		alu_inputs[6:1],
		alu_inputs[70:7] };
      default: IF_IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_ETC___d388 =
		   { 2'd3,
		     s3system_rs1_imm__h7842,
		     rx_stage1_control_first_x_BITS_63_TO_0__q5[1:0],
		     ff_stage1_meta_w_datawget_BITS_40_TO_9__q4[11:0],
		     ff_stage1_meta_w_datawget_BITS_8_TO_2__q3[2:0] };
    endcase
  end
  always@(ff_stage3_type_w_data_wget)
  begin
    case (ff_stage3_type_w_data_wget[67:66])
      2'd0, 2'd1:
	  IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435 =
	      ff_stage3_type_w_data_wget[67:66];
      2'd2: IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435 = 2'd3;
      2'd3: IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435 = 2'd2;
    endcase
  end
  always@(IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435)
  begin
    case (IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435)
      2'd0, 2'd1:
	  CASE_IF_ff_stage3_type_w_data_whas__23_THEN_IF_ETC__q6 =
	      IF_ff_stage3_type_w_data_whas__23_THEN_IF_ff_s_ETC___d435;
      2'd2: CASE_IF_ff_stage3_type_w_data_whas__23_THEN_IF_ETC__q6 = 2'd3;
      2'd3: CASE_IF_ff_stage3_type_w_data_whas__23_THEN_IF_ETC__q6 = 2'd2;
    endcase
  end
  always@(v_trigger_data1_1_wget)
  begin
    case (v_trigger_data1_1_wget[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_v_trigger_data1_1wget_BITS_21_TO_20_0_v__ETC__q7 =
	      v_trigger_data1_1_wget;
      2'd3:
	  CASE_v_trigger_data1_1wget_BITS_21_TO_20_0_v__ETC__q7 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(v_trigger_data1_0_wget)
  begin
    case (v_trigger_data1_0_wget[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_v_trigger_data1_0wget_BITS_21_TO_20_0_v__ETC__q8 =
	      v_trigger_data1_0_wget;
      2'd3:
	  CASE_v_trigger_data1_0wget_BITS_21_TO_20_0_v__ETC__q8 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_eEpoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_loadreserved_addr <= `BSV_ASSIGNMENT_DELAY
	    { 1'd0, 32'hAAAAAAAA /* unspecified value */  };
	rg_wEpoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_eEpoch_EN) rg_eEpoch <= `BSV_ASSIGNMENT_DELAY rg_eEpoch_D_IN;
	if (rg_loadreserved_addr_EN)
	  rg_loadreserved_addr <= `BSV_ASSIGNMENT_DELAY
	      rg_loadreserved_addr_D_IN;
	if (rg_wEpoch_EN) rg_wEpoch <= `BSV_ASSIGNMENT_DELAY rg_wEpoch_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_eEpoch = 1'h0;
    rg_loadreserved_addr = 33'h0AAAAAAAA;
    rg_wEpoch = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d30 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d31 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d32 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h3163 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("[%10d", v__h3163, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("STAGE2 : ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("TraceDump { ", "pc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("'h%h", rx_stage1_dump_first_x[95:32]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write(", ", "instruction: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("'h%h", rx_stage1_dump_first_x[31:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d30 ||
	   TASK_testplusargs___d31 && TASK_testplusargs___d32))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d42 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d43 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d44 = $test$plusargs("l1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h3348 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("[%10d", v__h3348, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("STAGE2 : OPs: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("STAGE1_operands { ", "op1: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("'h%h", rx_stage1_operands_first_x[127:64]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write(", ", "op2: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("'h%h", rx_stage1_operands_first_x[63:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d42 ||
	   TASK_testplusargs___d43 && TASK_testplusargs___d44))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d54 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d55 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d56 = $test$plusargs("l1");
	  #0;
	end
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d65 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd0;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d67 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd1;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d69 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd2;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d71 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd3;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d73 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd4;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d75 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd5;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d77 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd6;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d79 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd7;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d107 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 == 2'd1;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d95 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd0 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd1 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd2 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd3 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd4 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd5 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd6 &&
	ff_stage1_meta_w_data_wget[46:43] != 4'd7;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d105 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 == 2'd0;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d109 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 == 2'd2;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d115 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 != 2'd0 &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 != 2'd1 &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 != 2'd2;
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d123 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	!ff_stage1_meta_w_data_wget[1];
    TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d125 =
	(TASK_testplusargs___d54 ||
	 TASK_testplusargs___d55 && TASK_testplusargs___d56) &&
	ff_stage1_meta_w_data_wget[1];
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h3537 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("[%10d", v__h3537, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("STAGE2 : Meta: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("InstrMeta { ", "inst_type: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d65)
	$write("ALU");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d67)
	$write("MEMORY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d69)
	$write("BRANCH");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d71)
	$write("JAL");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d73)
	$write("JALR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d75)
	$write("SYSTEM_INSTR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d77)
	$write("TRAP");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d79)
	$write("WFI");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d95)
	$write("MULDIV");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write(", ", "memaccess: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d105)
	$write("Load");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d107)
	$write("Store");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d109)
	$write("Fence");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d115)
	$write("Atomic");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write(", ", "immediate: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("'h%h", ff_stage1_meta_w_data_wget[40:9]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write(", ", "funct: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("'h%h", ff_stage1_meta_w_data_wget[8:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write(", ", "word32: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d123)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_4_OR_TASK_testplusargs_5_AND_ETC___d125)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write(" }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d54 ||
	   TASK_testplusargs___d55 && TASK_testplusargs___d56))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d126 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d127 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d128 = $test$plusargs("l1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h3898 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("[%10d", v__h3898, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("STAGE2 : OpAddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("OpAddr { ", "rs1addr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("'h%h", ff_stage1_meta_w_data_wget[64:60]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write(", ", "rs2addr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("'h%h", ff_stage1_meta_w_data_wget[59:55]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write(", ", "rd: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("'h%h", ff_stage1_meta_w_data_wget[54:50], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d126 ||
	   TASK_testplusargs___d127 && TASK_testplusargs___d128))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d138 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d139 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d140 = $test$plusargs("l1");
	  #0;
	end
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d147 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	!ff_stage1_meta_w_data_wget[49];
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d149 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	ff_stage1_meta_w_data_wget[49];
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d153 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	ff_stage1_meta_w_data_wget[48:47] == 2'd0;
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d155 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	ff_stage1_meta_w_data_wget[48:47] == 2'd1;
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d157 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	ff_stage1_meta_w_data_wget[48:47] == 2'd2;
    TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d163 =
	(TASK_testplusargs___d138 ||
	 TASK_testplusargs___d139 && TASK_testplusargs___d140) &&
	ff_stage1_meta_w_data_wget[48:47] != 2'd0 &&
	ff_stage1_meta_w_data_wget[48:47] != 2'd1 &&
	ff_stage1_meta_w_data_wget[48:47] != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h4078 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write("[%10d", v__h4078, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write("STAGE2 : OpType: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write("OpType { ", "rs1type: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d147)
	$write("IntegerRF");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d149)
	$write("PC");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write(", ", "rs2type: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d153)
	$write("IntegerRF");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d155)
	$write("Immediate");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d157)
	$write("Constant4");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_38_OR_TASK_testplusargs_39_A_ETC___d163)
	$write("Constant2");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write(" }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d138 ||
	   TASK_testplusargs___d139 && TASK_testplusargs___d140))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d164 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d165 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d166 = $test$plusargs("l1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h4298 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("[%10d", v__h4298, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("STAGE2 : Control: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("STAGE1_control { ", "epoch: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("'h%h", rx_stage1_control_first_x[65:64]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write(", ", "pc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("'h%h", rx_stage1_control_first_x[63:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d164 ||
	   TASK_testplusargs___d165 && TASK_testplusargs___d166))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d176 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d177 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d178 = $test$plusargs("l1");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h4485 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d176 ||
	   TASK_testplusargs___d177 && TASK_testplusargs___d178))
	$write("[%10d", v__h4485, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d176 ||
	   TASK_testplusargs___d177 && TASK_testplusargs___d178))
	$write("STAGE2 : Fwding : Valid:%b Op1:%h Op2:%h",
	       NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195,
	       op1__h3084,
	       op2__h3085);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d176 ||
	   TASK_testplusargs___d177 && TASK_testplusargs___d178))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d239 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d240 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  TASK_testplusargs___d241 = $test$plusargs("l1");
	  #0;
	end
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d247 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[137];
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d249 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	!alu_inputs[137];
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d252 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[136:135] == 2'd0;
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d254 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[136:135] == 2'd1;
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d256 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[136:135] == 2'd2;
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d262 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[136:135] != 2'd0 &&
	alu_inputs[136:135] != 2'd1 &&
	alu_inputs[136:135] != 2'd2;
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d267 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	alu_inputs[0];
    TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d269 =
	(TASK_testplusargs___d239 ||
	 TASK_testplusargs___d240 && TASK_testplusargs___d241) &&
	!alu_inputs[0];
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass)
	begin
	  v__h6283 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("[%10d", v__h6283, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("STAGE2 : AluOut: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("ALU_OUT { ", "done: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d247)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d249)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(", ", "cmtype: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d252)
	$write("MEMORY");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d254)
	$write("SYSTEM_INSTR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d256)
	$write("REGULAR");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d262)
	$write("TRAP");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(", ", "aluresult: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("'h%h", alu_inputs[134:71]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(", ", "effective_addr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("'h%h", alu_inputs[70:7]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(", ", "cause: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("'h%h", alu_inputs[6:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(", ", "redirect: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d267)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  TASK_testplusargs_39_OR_TASK_testplusargs_40_A_ETC___d269)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write(" }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  (TASK_testplusargs___d239 ||
	   TASK_testplusargs___d240 && TASK_testplusargs___d241))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292)
	begin
	  TASK_testplusargs___d294 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292)
	begin
	  TASK_testplusargs___d295 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292)
	begin
	  TASK_testplusargs___d296 = $test$plusargs("l1");
	  #0;
	end
    IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d299 =
	x__h6827 == 5'b00101 &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_IF_ff_st_ETC___d103 == 2'd3 &&
	(TASK_testplusargs___d294 ||
	 TASK_testplusargs___d295 && TASK_testplusargs___d296);
    IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d302 =
	IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d299;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d292)
	begin
	  v__h6977 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d302)
	$write("[%10d", v__h6977, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d302)
	$write("STAGE2: Reserving Addr: %h", alu_inputs[70:7]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d302)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309)
	begin
	  TASK_testplusargs___d311 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309)
	begin
	  TASK_testplusargs___d312 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309)
	begin
	  TASK_testplusargs___d313 = $test$plusargs("l1");
	  #0;
	end
    IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d316 =
	x__h6827 == 5'b00111 &&
	IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 == 2'd3 &&
	(TASK_testplusargs___d311 ||
	 TASK_testplusargs___d312 && TASK_testplusargs___d313);
    TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d323 =
	(TASK_testplusargs___d311 ||
	 TASK_testplusargs___d312 && TASK_testplusargs___d313) &&
	rg_loadreserved_addr[32];
    TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d330 =
	(TASK_testplusargs___d311 ||
	 TASK_testplusargs___d312 && TASK_testplusargs___d313) &&
	!rg_loadreserved_addr[32];
    IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d319 =
	IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	IF_ff_stage1_meta_w_data_whas__0_THEN_ff_stage_ETC___d316;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d309)
	begin
	  v__h7230 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d319)
	$write("[%10d", v__h7230, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d319)
	$write("STAGE2: SC-ADDR:%h RES-ADDR: ", alu_inputs[70:7]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	  ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	  x__h6827 == 5'b00111 &&
	  IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 == 2'd3 &&
	  TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d323)
	$write("tagged Valid ", "'h%h", rg_loadreserved_addr[31:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	  NOT_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_s_ETC___d195 &&
	  ff_stage1_meta_w_data_wget[46:43] == 4'd1 &&
	  x__h6827 == 5'b00111 &&
	  IF_IF_ff_stage1_meta_w_data_whas__0_THEN_ff_st_ETC___d305 == 2'd3 &&
	  TASK_testplusargs_11_OR_TASK_testplusargs_12_A_ETC___d330)
	$write("tagged Invalid ", "");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d319)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  !IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273)
	begin
	  TASK_testplusargs___d391 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  !IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273)
	begin
	  TASK_testplusargs___d392 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  !IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273)
	begin
	  TASK_testplusargs___d393 = $test$plusargs("l0");
	  #0;
	end
    NOT_IF_ff_stage1_control_w_data_whas__70_THEN__ETC___d396 =
	!IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273 &&
	(TASK_testplusargs___d391 ||
	 TASK_testplusargs___d392 && TASK_testplusargs___d393);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  !IF_ff_stage1_control_w_data_whas__70_THEN_ff_s_ETC___d273)
	begin
	  v__h6617 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  NOT_IF_ff_stage1_control_w_data_whas__70_THEN__ETC___d396)
	$write("[%10d", v__h6617, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  NOT_IF_ff_stage1_control_w_data_whas__70_THEN__ETC___d396)
	$write("STAGE2 : Dropping instruction due to mis - match");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_fetch_execute_pass &&
	  NOT_IF_ff_stage1_control_w_data_whas__70_THEN__ETC___d396)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch)
	begin
	  TASK_testplusargs___d470 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch)
	begin
	  TASK_testplusargs___d471 = $test$plusargs("mstage2");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch)
	begin
	  TASK_testplusargs___d472 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch)
	begin
	  v__h9106 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch &&
	  (TASK_testplusargs___d470 ||
	   TASK_testplusargs___d471 && TASK_testplusargs___d472))
	$write("[%10d", v__h9106, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch &&
	  (TASK_testplusargs___d470 ||
	   TASK_testplusargs___d471 && TASK_testplusargs___d472))
	$write("STAGE2: Received Flush from WB");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_ma_update_wEpoch &&
	  (TASK_testplusargs___d470 ||
	   TASK_testplusargs___d471 && TASK_testplusargs___d472))
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkstage2

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:11 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// rx_stage3_common_deq_ena       O     1
// rx_stage3_type_deq_ena         O     1
// rx_stage3_dump_deq_ena         O     1
// RDY_memory_response_put        O     1 const
// commit_rd_get                  O    69
// RDY_commit_rd_get              O     1
// operand_fwding_get             O    70
// RDY_operand_fwding_get         O     1 const
// flush_fst                      O    64
// RDY_flush_fst                  O     1 const
// flush_snd                      O     1
// RDY_flush_snd                  O     1 const
// mv_csr_decode                  O   152
// RDY_mv_csr_decode              O     1 const
// mv_csr_misa_c                  O     1 reg
// RDY_mv_csr_misa_c              O     1 const
// RDY_clint_msip                 O     1 const
// RDY_clint_mtip                 O     1 const
// RDY_clint_mtime                O     1 const
// RDY_ext_interrupt              O     1 const
// csr_updated                    O     1 const
// RDY_csr_updated                O     1 const
// mv_interrupt                   O     1
// dump_get                       O   167
// RDY_dump_get                   O     1 reg
// mv_trigger_data1               O    44
// RDY_mv_trigger_data1           O     1 const
// mv_trigger_data2               O   128 reg
// RDY_mv_trigger_data2           O     1 const
// mv_trigger_enable              O     2
// RDY_mv_trigger_enable          O     1 const
// mv_curr_priv                   O     2
// RDY_mv_curr_priv               O     1 const
// RDY_ma_delayed_output          O     1 const
// mv_pmp_cfg                     O    32 reg
// RDY_mv_pmp_cfg                 O     1 const
// mv_pmp_addr                    O   120 reg
// RDY_mv_pmp_addr                O     1 const
// CLK                            I     1 clock
// RST_N                          I     1 reset
// rx_stage3_common_notEmpty_b    I     1 unused
// rx_stage3_common_first_deq_rdy_b  I     1
// rx_stage3_common_first_x       I    70
// rx_stage3_type_notEmpty_b      I     1 unused
// rx_stage3_type_first_deq_rdy_b  I     1
// rx_stage3_type_first_x         I    83
// rx_stage3_dump_notEmpty_b      I     1 unused
// rx_stage3_dump_first_deq_rdy_b  I     1
// rx_stage3_dump_first_x         I    96
// memory_response_put            I    66
// clint_msip_intrpt              I     1 reg
// clint_mtip_intrpt              I     1 reg
// clint_mtime_c_mtime            I    64 reg
// ext_interrupt_i                I     1 reg
// ma_delayed_output_r            I    65
// EN_memory_response_put         I     1
// EN_clint_msip                  I     1
// EN_clint_mtip                  I     1
// EN_clint_mtime                 I     1
// EN_ext_interrupt               I     1
// EN_ma_delayed_output           I     1
// EN_commit_rd_get               I     1 unused
// EN_operand_fwding_get          I     1 unused
// EN_dump_get                    I     1
//
// Combinational paths from inputs to outputs:
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> rx_stage3_common_deq_ena
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> rx_stage3_type_deq_ena
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> rx_stage3_dump_deq_ena
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> RDY_commit_rd_get
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    EN_ma_delayed_output,
//    EN_dump_get) -> flush_fst
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    EN_ma_delayed_output,
//    EN_dump_get) -> flush_snd
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> commit_rd_get
//   (rx_stage3_common_first_deq_rdy_b,
//    rx_stage3_common_first_x,
//    rx_stage3_type_first_deq_rdy_b,
//    rx_stage3_type_first_x,
//    rx_stage3_dump_first_deq_rdy_b,
//    ma_delayed_output_r,
//    EN_ma_delayed_output,
//    EN_dump_get) -> operand_fwding_get
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkstage3(CLK,
		RST_N,

		rx_stage3_common_notEmpty_b,

		rx_stage3_common_first_deq_rdy_b,

		rx_stage3_common_first_x,

		rx_stage3_common_deq_ena,

		rx_stage3_type_notEmpty_b,

		rx_stage3_type_first_deq_rdy_b,

		rx_stage3_type_first_x,

		rx_stage3_type_deq_ena,

		rx_stage3_dump_notEmpty_b,

		rx_stage3_dump_first_deq_rdy_b,

		rx_stage3_dump_first_x,

		rx_stage3_dump_deq_ena,

		memory_response_put,
		EN_memory_response_put,
		RDY_memory_response_put,

		EN_commit_rd_get,
		commit_rd_get,
		RDY_commit_rd_get,

		EN_operand_fwding_get,
		operand_fwding_get,
		RDY_operand_fwding_get,

		flush_fst,
		RDY_flush_fst,

		flush_snd,
		RDY_flush_snd,

		mv_csr_decode,
		RDY_mv_csr_decode,

		mv_csr_misa_c,
		RDY_mv_csr_misa_c,

		clint_msip_intrpt,
		EN_clint_msip,
		RDY_clint_msip,

		clint_mtip_intrpt,
		EN_clint_mtip,
		RDY_clint_mtip,

		clint_mtime_c_mtime,
		EN_clint_mtime,
		RDY_clint_mtime,

		ext_interrupt_i,
		EN_ext_interrupt,
		RDY_ext_interrupt,

		csr_updated,
		RDY_csr_updated,

		mv_interrupt,

		EN_dump_get,
		dump_get,
		RDY_dump_get,

		mv_trigger_data1,
		RDY_mv_trigger_data1,

		mv_trigger_data2,
		RDY_mv_trigger_data2,

		mv_trigger_enable,
		RDY_mv_trigger_enable,

		mv_curr_priv,
		RDY_mv_curr_priv,

		ma_delayed_output_r,
		EN_ma_delayed_output,
		RDY_ma_delayed_output,

		mv_pmp_cfg,
		RDY_mv_pmp_cfg,

		mv_pmp_addr,
		RDY_mv_pmp_addr);
  input  CLK;
  input  RST_N;

  // action method rx_stage3_common_notEmpty
  input  rx_stage3_common_notEmpty_b;

  // action method rx_stage3_common_first_deq_rdy
  input  rx_stage3_common_first_deq_rdy_b;

  // action method rx_stage3_common_first
  input  [69 : 0] rx_stage3_common_first_x;

  // value method rx_stage3_common_deq_ena
  output rx_stage3_common_deq_ena;

  // action method rx_stage3_type_notEmpty
  input  rx_stage3_type_notEmpty_b;

  // action method rx_stage3_type_first_deq_rdy
  input  rx_stage3_type_first_deq_rdy_b;

  // action method rx_stage3_type_first
  input  [82 : 0] rx_stage3_type_first_x;

  // value method rx_stage3_type_deq_ena
  output rx_stage3_type_deq_ena;

  // action method rx_stage3_dump_notEmpty
  input  rx_stage3_dump_notEmpty_b;

  // action method rx_stage3_dump_first_deq_rdy
  input  rx_stage3_dump_first_deq_rdy_b;

  // action method rx_stage3_dump_first
  input  [95 : 0] rx_stage3_dump_first_x;

  // value method rx_stage3_dump_deq_ena
  output rx_stage3_dump_deq_ena;

  // action method memory_response_put
  input  [65 : 0] memory_response_put;
  input  EN_memory_response_put;
  output RDY_memory_response_put;

  // actionvalue method commit_rd_get
  input  EN_commit_rd_get;
  output [68 : 0] commit_rd_get;
  output RDY_commit_rd_get;

  // actionvalue method operand_fwding_get
  input  EN_operand_fwding_get;
  output [69 : 0] operand_fwding_get;
  output RDY_operand_fwding_get;

  // value method flush_fst
  output [63 : 0] flush_fst;
  output RDY_flush_fst;

  // value method flush_snd
  output flush_snd;
  output RDY_flush_snd;

  // value method mv_csr_decode
  output [151 : 0] mv_csr_decode;
  output RDY_mv_csr_decode;

  // value method mv_csr_misa_c
  output mv_csr_misa_c;
  output RDY_mv_csr_misa_c;

  // action method clint_msip
  input  clint_msip_intrpt;
  input  EN_clint_msip;
  output RDY_clint_msip;

  // action method clint_mtip
  input  clint_mtip_intrpt;
  input  EN_clint_mtip;
  output RDY_clint_mtip;

  // action method clint_mtime
  input  [63 : 0] clint_mtime_c_mtime;
  input  EN_clint_mtime;
  output RDY_clint_mtime;

  // action method ext_interrupt
  input  ext_interrupt_i;
  input  EN_ext_interrupt;
  output RDY_ext_interrupt;

  // value method csr_updated
  output csr_updated;
  output RDY_csr_updated;

  // value method mv_interrupt
  output mv_interrupt;

  // actionvalue method dump_get
  input  EN_dump_get;
  output [166 : 0] dump_get;
  output RDY_dump_get;

  // value method mv_trigger_data1
  output [43 : 0] mv_trigger_data1;
  output RDY_mv_trigger_data1;

  // value method mv_trigger_data2
  output [127 : 0] mv_trigger_data2;
  output RDY_mv_trigger_data2;

  // value method mv_trigger_enable
  output [1 : 0] mv_trigger_enable;
  output RDY_mv_trigger_enable;

  // value method mv_curr_priv
  output [1 : 0] mv_curr_priv;
  output RDY_mv_curr_priv;

  // action method ma_delayed_output
  input  [64 : 0] ma_delayed_output_r;
  input  EN_ma_delayed_output;
  output RDY_ma_delayed_output;

  // value method mv_pmp_cfg
  output [31 : 0] mv_pmp_cfg;
  output RDY_mv_pmp_cfg;

  // value method mv_pmp_addr
  output [119 : 0] mv_pmp_addr;
  output RDY_mv_pmp_addr;

  // signals for module outputs
  wire [166 : 0] dump_get;
  wire [151 : 0] mv_csr_decode;
  wire [127 : 0] mv_trigger_data2;
  wire [119 : 0] mv_pmp_addr;
  wire [69 : 0] operand_fwding_get;
  wire [68 : 0] commit_rd_get;
  wire [63 : 0] flush_fst;
  wire [43 : 0] mv_trigger_data1;
  wire [31 : 0] mv_pmp_cfg;
  wire [1 : 0] mv_curr_priv, mv_trigger_enable;
  wire RDY_clint_msip,
       RDY_clint_mtime,
       RDY_clint_mtip,
       RDY_commit_rd_get,
       RDY_csr_updated,
       RDY_dump_get,
       RDY_ext_interrupt,
       RDY_flush_fst,
       RDY_flush_snd,
       RDY_ma_delayed_output,
       RDY_memory_response_put,
       RDY_mv_csr_decode,
       RDY_mv_csr_misa_c,
       RDY_mv_curr_priv,
       RDY_mv_pmp_addr,
       RDY_mv_pmp_cfg,
       RDY_mv_trigger_data1,
       RDY_mv_trigger_data2,
       RDY_mv_trigger_enable,
       RDY_operand_fwding_get,
       csr_updated,
       flush_snd,
       mv_csr_misa_c,
       mv_interrupt,
       rx_stage3_common_deq_ena,
       rx_stage3_dump_deq_ena,
       rx_stage3_type_deq_ena;

  // inlined wires
  wire [82 : 0] ff_stage3_type_w_data_wget;
  wire [69 : 0] wr_commit_wget, wr_operand_fwding_wget;
  wire [66 : 0] wr_memory_response_1_wget;
  wire [64 : 0] wr_flush_wget;
  wire ff_stage3_common_w_ena_whas,
       ff_stage3_dump_w_ena_whas,
       ff_stage3_type_w_ena_whas,
       wr_commit_whas,
       wr_flush_whas,
       wr_operand_fwding_whas;

  // register rg_epoch
  reg rg_epoch;
  wire rg_epoch_D_IN, rg_epoch_EN;

  // register rg_rerun
  reg rg_rerun;
  wire rg_rerun_D_IN, rg_rerun_EN;

  // register wr_memory_response
  reg [66 : 0] wr_memory_response;
  wire [66 : 0] wr_memory_response_D_IN;
  wire wr_memory_response_EN;

  // ports of submodule csr
  wire [151 : 0] csr_mv_csr_decode;
  wire [128 : 0] csr_system_instruction;
  wire [127 : 0] csr_mv_trigger_data2;
  wire [119 : 0] csr_mv_pmp_addr;
  wire [63 : 0] csr_clint_mtime_c_mtime,
		csr_system_instruction_op1,
		csr_take_trap,
		csr_take_trap_badaddr,
		csr_take_trap_pc;
  wire [43 : 0] csr_mv_trigger_data1;
  wire [31 : 0] csr_mv_pmp_cfg;
  wire [11 : 0] csr_system_instruction_csr_address;
  wire [5 : 0] csr_take_trap_type_cause;
  wire [2 : 0] csr_system_instruction_funct3;
  wire [1 : 0] csr_mv_curr_priv,
	       csr_mv_trigger_enable,
	       csr_system_instruction_lpc;
  wire csr_EN_clint_msip,
       csr_EN_clint_mtime,
       csr_EN_clint_mtip,
       csr_EN_ext_interrupt,
       csr_EN_incr_minstret,
       csr_EN_system_instruction,
       csr_EN_take_trap,
       csr_clint_msip_intrpt,
       csr_clint_mtip_intrpt,
       csr_ext_interrupt_ex_i,
       csr_mv_csr_misa_c,
       csr_mv_interrupt;

  // ports of submodule dump_ff
  wire [166 : 0] dump_ff_D_IN, dump_ff_D_OUT;
  wire dump_ff_CLR, dump_ff_DEQ, dump_ff_EMPTY_N, dump_ff_ENQ, dump_ff_FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_increment_instruction_counter,
       CAN_FIRE_RL_instruction_commit,
       CAN_FIRE_RL_wr_memory_response__dreg_update,
       CAN_FIRE_clint_msip,
       CAN_FIRE_clint_mtime,
       CAN_FIRE_clint_mtip,
       CAN_FIRE_commit_rd_get,
       CAN_FIRE_dump_get,
       CAN_FIRE_ext_interrupt,
       CAN_FIRE_ma_delayed_output,
       CAN_FIRE_memory_response_put,
       CAN_FIRE_operand_fwding_get,
       CAN_FIRE_rx_stage3_common_first,
       CAN_FIRE_rx_stage3_common_first_deq_rdy,
       CAN_FIRE_rx_stage3_common_notEmpty,
       CAN_FIRE_rx_stage3_dump_first,
       CAN_FIRE_rx_stage3_dump_first_deq_rdy,
       CAN_FIRE_rx_stage3_dump_notEmpty,
       CAN_FIRE_rx_stage3_type_first,
       CAN_FIRE_rx_stage3_type_first_deq_rdy,
       CAN_FIRE_rx_stage3_type_notEmpty,
       WILL_FIRE_RL_increment_instruction_counter,
       WILL_FIRE_RL_instruction_commit,
       WILL_FIRE_RL_wr_memory_response__dreg_update,
       WILL_FIRE_clint_msip,
       WILL_FIRE_clint_mtime,
       WILL_FIRE_clint_mtip,
       WILL_FIRE_commit_rd_get,
       WILL_FIRE_dump_get,
       WILL_FIRE_ext_interrupt,
       WILL_FIRE_ma_delayed_output,
       WILL_FIRE_memory_response_put,
       WILL_FIRE_operand_fwding_get,
       WILL_FIRE_rx_stage3_common_first,
       WILL_FIRE_rx_stage3_common_first_deq_rdy,
       WILL_FIRE_rx_stage3_common_notEmpty,
       WILL_FIRE_rx_stage3_dump_first,
       WILL_FIRE_rx_stage3_dump_first_deq_rdy,
       WILL_FIRE_rx_stage3_dump_notEmpty,
       WILL_FIRE_rx_stage3_type_first,
       WILL_FIRE_rx_stage3_type_first_deq_rdy,
       WILL_FIRE_rx_stage3_type_notEmpty;

  // declarations used by system tasks
  // synopsys translate_off
  reg TASK_testplusargs___d19;
  reg TASK_testplusargs___d20;
  reg TASK_testplusargs___d21;
  reg [63 : 0] v__h1870;
  reg TASK_testplusargs___d31;
  reg TASK_testplusargs___d32;
  reg TASK_testplusargs___d33;
  reg [63 : 0] v__h2055;
  reg TASK_testplusargs___d45;
  reg TASK_testplusargs___d46;
  reg TASK_testplusargs___d47;
  reg [63 : 0] v__h2250;
  reg TASK_testplusargs___d144;
  reg TASK_testplusargs___d145;
  reg TASK_testplusargs___d146;
  reg [63 : 0] v__h3248;
  reg TASK_testplusargs___d154;
  reg TASK_testplusargs___d155;
  reg TASK_testplusargs___d156;
  reg [63 : 0] v__h2907;
  reg TASK_testplusargs___d192;
  reg TASK_testplusargs___d193;
  reg TASK_testplusargs___d194;
  reg [63 : 0] v__h3730;
  reg TASK_testplusargs___d248;
  reg TASK_testplusargs___d249;
  reg TASK_testplusargs___d250;
  reg [63 : 0] v__h4969;
  reg TASK_testplusargs___d272;
  reg TASK_testplusargs___d273;
  reg TASK_testplusargs___d274;
  reg [63 : 0] v__h5043;
  reg TASK_testplusargs___d283;
  reg TASK_testplusargs___d284;
  reg TASK_testplusargs___d285;
  reg [63 : 0] v__h5138;
  reg rg_rerun_22_AND_TASK_testplusargs_44_OR_TASK_t_ETC___d149;
  reg ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d159;
  reg ff_stage3_type_w_data_wget__2_BIT_0_3_AND_NOT__ETC___d197;
  reg NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d199;
  reg wr_memory_response_15_BIT_1_20_AND_TASK_testpl_ETC___d253;
  reg NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d257;
  reg NOT_wr_memory_response_15_BIT_66_16_65_OR_NOT__ETC___d277;
  reg NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d280;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d85;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d88;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d106;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d109;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d112;
  reg TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d119;
  reg NOT_rg_epoch_24_EQ_IF_ff_stage3_common_w_data__ETC___d288;
  // synopsys translate_on

  // remaining internal signals
  reg [21 : 0] CASE_csrmv_trigger_data1_BITS_21_TO_20_0_csr_ETC__q2,
	       CASE_csrmv_trigger_data1_BITS_43_TO_42_0_csr_ETC__q1;
  reg [1 : 0] CASE_rx_stage3_type_first_x_BITS_67_TO_66_0_rx_ETC__q4,
	      CASE_rx_stage3_type_first_x_BITS_82_TO_81_0_rx_ETC__q3,
	      IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103;
  wire [166 : 0] _dfoo2;
  wire [100 : 0] IF_ff_stage3_dump_w_data_whas__5_THEN_ff_stage_ETC___d237;
  wire [69 : 0] _dfoo10;
  wire [64 : 0] _dfoo14;
  wire [63 : 0] _theResult_____1_snd__h3364,
		_theResult____h3307,
		_theResult____h4120,
		_theResult____h4431,
		data__h3311,
		x__read_rdvalue__h5759;
  wire [5 : 0] type_cause__h4513;
  wire [4 : 0] x__read_rdaddr__h5758;
  wire [1 : 0] IF_csr_mv_curr_priv__83_EQ_3_84_THEN_csr_mv_cu_ETC___d185;
  wire NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179,
       NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190,
       NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202,
       _dfoo1,
       _dfoo25,
       _dfoo3,
       _dfoo31,
       _dfoo33,
       _dfoo37,
       _dfoo39,
       _dfoo41,
       ff_stage3_type_w_data_whas__1_AND_NOT_ff_stage_ETC___d204,
       ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d224,
       ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d233,
       ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243,
       ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269,
       rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125,
       rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d128,
       rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153,
       rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d164,
       rg_rerun_22_OR_ff_stage3_type_w_data_whas__1_A_ETC___d127,
       wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218,
       x__h4837;

  // action method rx_stage3_common_notEmpty
  assign CAN_FIRE_rx_stage3_common_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage3_common_notEmpty = 1'd1 ;

  // action method rx_stage3_common_first_deq_rdy
  assign CAN_FIRE_rx_stage3_common_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage3_common_first_deq_rdy = 1'd1 ;

  // action method rx_stage3_common_first
  assign CAN_FIRE_rx_stage3_common_first = 1'd1 ;
  assign WILL_FIRE_rx_stage3_common_first = 1'd1 ;

  // value method rx_stage3_common_deq_ena
  assign rx_stage3_common_deq_ena = ff_stage3_common_w_ena_whas ;

  // action method rx_stage3_type_notEmpty
  assign CAN_FIRE_rx_stage3_type_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage3_type_notEmpty = 1'd1 ;

  // action method rx_stage3_type_first_deq_rdy
  assign CAN_FIRE_rx_stage3_type_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage3_type_first_deq_rdy = 1'd1 ;

  // action method rx_stage3_type_first
  assign CAN_FIRE_rx_stage3_type_first = 1'd1 ;
  assign WILL_FIRE_rx_stage3_type_first = 1'd1 ;

  // value method rx_stage3_type_deq_ena
  assign rx_stage3_type_deq_ena = ff_stage3_type_w_ena_whas ;

  // action method rx_stage3_dump_notEmpty
  assign CAN_FIRE_rx_stage3_dump_notEmpty = 1'd1 ;
  assign WILL_FIRE_rx_stage3_dump_notEmpty = 1'd1 ;

  // action method rx_stage3_dump_first_deq_rdy
  assign CAN_FIRE_rx_stage3_dump_first_deq_rdy = 1'd1 ;
  assign WILL_FIRE_rx_stage3_dump_first_deq_rdy = 1'd1 ;

  // action method rx_stage3_dump_first
  assign CAN_FIRE_rx_stage3_dump_first = 1'd1 ;
  assign WILL_FIRE_rx_stage3_dump_first = 1'd1 ;

  // value method rx_stage3_dump_deq_ena
  assign rx_stage3_dump_deq_ena = ff_stage3_dump_w_ena_whas ;

  // action method memory_response_put
  assign RDY_memory_response_put = 1'd1 ;
  assign CAN_FIRE_memory_response_put = 1'd1 ;
  assign WILL_FIRE_memory_response_put = EN_memory_response_put ;

  // actionvalue method commit_rd_get
  assign commit_rd_get = wr_commit_wget[68:0] ;
  assign RDY_commit_rd_get = wr_commit_whas && wr_commit_wget[69] ;
  assign CAN_FIRE_commit_rd_get = RDY_commit_rd_get ;
  assign WILL_FIRE_commit_rd_get = EN_commit_rd_get ;

  // actionvalue method operand_fwding_get
  assign operand_fwding_get =
	     { x__read_rdaddr__h5758,
	       x__read_rdvalue__h5759,
	       wr_operand_fwding_whas && wr_operand_fwding_wget[0] } ;
  assign RDY_operand_fwding_get = 1'd1 ;
  assign CAN_FIRE_operand_fwding_get = 1'd1 ;
  assign WILL_FIRE_operand_fwding_get = EN_operand_fwding_get ;

  // value method flush_fst
  assign flush_fst = wr_flush_wget[64:1] ;
  assign RDY_flush_fst = 1'd1 ;

  // value method flush_snd
  assign flush_snd = wr_flush_whas && wr_flush_wget[0] ;
  assign RDY_flush_snd = 1'd1 ;

  // value method mv_csr_decode
  assign mv_csr_decode =
	     { (csr_mv_csr_decode[151:150] == 2'd3) ?
		 csr_mv_csr_decode[151:150] :
		 2'd0,
	       csr_mv_csr_decode[149:0] } ;
  assign RDY_mv_csr_decode = 1'd1 ;

  // value method mv_csr_misa_c
  assign mv_csr_misa_c = csr_mv_csr_misa_c ;
  assign RDY_mv_csr_misa_c = 1'd1 ;

  // action method clint_msip
  assign RDY_clint_msip = 1'd1 ;
  assign CAN_FIRE_clint_msip = 1'd1 ;
  assign WILL_FIRE_clint_msip = EN_clint_msip ;

  // action method clint_mtip
  assign RDY_clint_mtip = 1'd1 ;
  assign CAN_FIRE_clint_mtip = 1'd1 ;
  assign WILL_FIRE_clint_mtip = EN_clint_mtip ;

  // action method clint_mtime
  assign RDY_clint_mtime = 1'd1 ;
  assign CAN_FIRE_clint_mtime = 1'd1 ;
  assign WILL_FIRE_clint_mtime = EN_clint_mtime ;

  // action method ext_interrupt
  assign RDY_ext_interrupt = 1'd1 ;
  assign CAN_FIRE_ext_interrupt = 1'd1 ;
  assign WILL_FIRE_ext_interrupt = EN_ext_interrupt ;

  // value method csr_updated
  assign csr_updated = 1'b0 ;
  assign RDY_csr_updated = 1'd1 ;

  // value method mv_interrupt
  assign mv_interrupt = csr_mv_interrupt ;

  // actionvalue method dump_get
  assign dump_get =
	     { (dump_ff_D_OUT[166:165] == 2'd3) ?
		 dump_ff_D_OUT[166:165] :
		 2'd0,
	       dump_ff_D_OUT[164:0] } ;
  assign RDY_dump_get = dump_ff_EMPTY_N ;
  assign CAN_FIRE_dump_get = dump_ff_EMPTY_N ;
  assign WILL_FIRE_dump_get = EN_dump_get ;

  // value method mv_trigger_data1
  assign mv_trigger_data1 =
	     { CASE_csrmv_trigger_data1_BITS_43_TO_42_0_csr_ETC__q1,
	       CASE_csrmv_trigger_data1_BITS_21_TO_20_0_csr_ETC__q2 } ;
  assign RDY_mv_trigger_data1 = 1'd1 ;

  // value method mv_trigger_data2
  assign mv_trigger_data2 = csr_mv_trigger_data2 ;
  assign RDY_mv_trigger_data2 = 1'd1 ;

  // value method mv_trigger_enable
  assign mv_trigger_enable = csr_mv_trigger_enable ;
  assign RDY_mv_trigger_enable = 1'd1 ;

  // value method mv_curr_priv
  assign mv_curr_priv = csr_mv_curr_priv ;
  assign RDY_mv_curr_priv = 1'd1 ;

  // action method ma_delayed_output
  assign RDY_ma_delayed_output = 1'd1 ;
  assign CAN_FIRE_ma_delayed_output = 1'd1 ;
  assign WILL_FIRE_ma_delayed_output = EN_ma_delayed_output ;

  // value method mv_pmp_cfg
  assign mv_pmp_cfg = csr_mv_pmp_cfg ;
  assign RDY_mv_pmp_cfg = 1'd1 ;

  // value method mv_pmp_addr
  assign mv_pmp_addr = csr_mv_pmp_addr ;
  assign RDY_mv_pmp_addr = 1'd1 ;

  // submodule csr
  mkcsr csr(.CLK(CLK),
	    .RST_N(RST_N),
	    .clint_msip_intrpt(csr_clint_msip_intrpt),
	    .clint_mtime_c_mtime(csr_clint_mtime_c_mtime),
	    .clint_mtip_intrpt(csr_clint_mtip_intrpt),
	    .ext_interrupt_ex_i(csr_ext_interrupt_ex_i),
	    .system_instruction_csr_address(csr_system_instruction_csr_address),
	    .system_instruction_funct3(csr_system_instruction_funct3),
	    .system_instruction_lpc(csr_system_instruction_lpc),
	    .system_instruction_op1(csr_system_instruction_op1),
	    .take_trap_badaddr(csr_take_trap_badaddr),
	    .take_trap_pc(csr_take_trap_pc),
	    .take_trap_type_cause(csr_take_trap_type_cause),
	    .EN_system_instruction(csr_EN_system_instruction),
	    .EN_take_trap(csr_EN_take_trap),
	    .EN_clint_msip(csr_EN_clint_msip),
	    .EN_clint_mtip(csr_EN_clint_mtip),
	    .EN_clint_mtime(csr_EN_clint_mtime),
	    .EN_incr_minstret(csr_EN_incr_minstret),
	    .EN_ext_interrupt(csr_EN_ext_interrupt),
	    .system_instruction(csr_system_instruction),
	    .RDY_system_instruction(),
	    .mv_csr_decode(csr_mv_csr_decode),
	    .RDY_mv_csr_decode(),
	    .take_trap(csr_take_trap),
	    .RDY_take_trap(),
	    .RDY_clint_msip(),
	    .RDY_clint_mtip(),
	    .RDY_clint_mtime(),
	    .RDY_incr_minstret(),
	    .RDY_ext_interrupt(),
	    .mv_csr_misa_c(csr_mv_csr_misa_c),
	    .RDY_mv_csr_misa_c(),
	    .mv_interrupt(csr_mv_interrupt),
	    .mv_curr_priv(csr_mv_curr_priv),
	    .RDY_mv_curr_priv(),
	    .csr_mstatus(),
	    .RDY_csr_mstatus(),
	    .mv_pmp_cfg(csr_mv_pmp_cfg),
	    .RDY_mv_pmp_cfg(),
	    .mv_pmp_addr(csr_mv_pmp_addr),
	    .RDY_mv_pmp_addr(),
	    .mv_trigger_data1(csr_mv_trigger_data1),
	    .RDY_mv_trigger_data1(),
	    .mv_trigger_data2(csr_mv_trigger_data2),
	    .RDY_mv_trigger_data2(),
	    .mv_trigger_enable(csr_mv_trigger_enable),
	    .RDY_mv_trigger_enable());

  // submodule dump_ff
  FIFOL1 #(.width(32'd167)) dump_ff(.RST(RST_N),
				    .CLK(CLK),
				    .D_IN(dump_ff_D_IN),
				    .ENQ(dump_ff_ENQ),
				    .DEQ(dump_ff_DEQ),
				    .CLR(dump_ff_CLR),
				    .D_OUT(dump_ff_D_OUT),
				    .FULL_N(dump_ff_FULL_N),
				    .EMPTY_N(dump_ff_EMPTY_N));

  // rule RL_instruction_commit
  assign CAN_FIRE_RL_instruction_commit =
	     rx_stage3_common_first_deq_rdy_b &&
	     rx_stage3_type_first_deq_rdy_b &&
	     rx_stage3_dump_first_deq_rdy_b &&
	     EN_ma_delayed_output &&
	     dump_ff_FULL_N ;
  assign WILL_FIRE_RL_instruction_commit = CAN_FIRE_RL_instruction_commit ;

  // rule RL_increment_instruction_counter
  assign CAN_FIRE_RL_increment_instruction_counter = RDY_commit_rd_get ;
  assign WILL_FIRE_RL_increment_instruction_counter =
	     CAN_FIRE_RL_increment_instruction_counter &&
	     !WILL_FIRE_RL_instruction_commit ;

  // rule RL_wr_memory_response__dreg_update
  assign CAN_FIRE_RL_wr_memory_response__dreg_update = 1'd1 ;
  assign WILL_FIRE_RL_wr_memory_response__dreg_update = 1'd1 ;

  // inlined wires
  assign ff_stage3_common_w_ena_whas =
	     WILL_FIRE_RL_instruction_commit && _dfoo41 ;
  assign ff_stage3_type_w_ena_whas =
	     WILL_FIRE_RL_instruction_commit && _dfoo39 ;
  assign ff_stage3_type_w_data_wget =
	     { CASE_rx_stage3_type_first_x_BITS_82_TO_81_0_rx_ETC__q3,
	       (rx_stage3_type_first_x[82:81] == 2'd0) ?
		 { 13'b0101010101010 /* unspecified value */ ,
		   CASE_rx_stage3_type_first_x_BITS_67_TO_66_0_rx_ETC__q4,
		   rx_stage3_type_first_x[65:0] } :
		 rx_stage3_type_first_x[80:0] } ;
  assign ff_stage3_dump_w_ena_whas =
	     WILL_FIRE_RL_instruction_commit && _dfoo37 ;
  assign wr_memory_response_1_wget = { 1'd1, memory_response_put } ;
  assign wr_operand_fwding_wget =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d164 ?
	       { rx_stage3_common_first_x[5:1],
		 data__h3311,
		 !ff_stage3_type_w_data_wget[0] || ma_delayed_output_r[0] } :
	       { rx_stage3_common_first_x[5:1], _theResult____h4431, 1'd1 } ;
  assign wr_operand_fwding_whas = WILL_FIRE_RL_instruction_commit && _dfoo25 ;
  assign wr_commit_wget =
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179) ?
	       { 1'd1, rx_stage3_common_first_x[5:1], data__h3311 } :
	       _dfoo10 ;
  assign wr_commit_whas =
	     WILL_FIRE_RL_instruction_commit &&
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 ||
	      _dfoo1) ;
  assign wr_flush_wget =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d128 ?
	       { rg_rerun ? rx_stage3_common_first_x[69:6] : csr_take_trap,
		 1'd1 } :
	       _dfoo14 ;
  assign wr_flush_whas = WILL_FIRE_RL_instruction_commit && _dfoo33 ;

  // register rg_epoch
  assign rg_epoch_D_IN = x__h4837 ;
  assign rg_epoch_EN = WILL_FIRE_RL_instruction_commit && _dfoo33 ;

  // register rg_rerun
  assign rg_rerun_D_IN =
	     !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 ||
	     !rg_rerun ;
  assign rg_rerun_EN = WILL_FIRE_RL_instruction_commit && _dfoo31 ;

  // register wr_memory_response
  assign wr_memory_response_D_IN =
	     { EN_memory_response_put && wr_memory_response_1_wget[66],
	       wr_memory_response_1_wget[65:0] } ;
  assign wr_memory_response_EN = 1'd1 ;

  // submodule csr
  assign csr_clint_msip_intrpt = clint_msip_intrpt ;
  assign csr_clint_mtime_c_mtime = clint_mtime_c_mtime ;
  assign csr_clint_mtip_intrpt = clint_mtip_intrpt ;
  assign csr_ext_interrupt_ex_i = ext_interrupt_i ;
  assign csr_system_instruction_csr_address =
	     ff_stage3_type_w_data_wget[14:3] ;
  assign csr_system_instruction_funct3 = ff_stage3_type_w_data_wget[2:0] ;
  assign csr_system_instruction_lpc = ff_stage3_type_w_data_wget[16:15] ;
  assign csr_system_instruction_op1 = ff_stage3_type_w_data_wget[80:17] ;
  assign csr_take_trap_badaddr =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153 ?
	       ff_stage3_type_w_data_wget[63:0] :
	       wr_memory_response[65:2] ;
  assign csr_take_trap_pc = rx_stage3_common_first_x[69:6] ;
  assign csr_take_trap_type_cause =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153 ?
	       ff_stage3_type_w_data_wget[69:64] :
	       type_cause__h4513 ;
  assign csr_EN_system_instruction =
	     WILL_FIRE_RL_instruction_commit &&
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202 ;
  assign csr_EN_take_trap =
	     WILL_FIRE_RL_instruction_commit &&
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153 ||
	      rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      !rg_rerun &&
	      ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243) ;
  assign csr_EN_clint_msip = EN_clint_msip ;
  assign csr_EN_clint_mtip = EN_clint_mtip ;
  assign csr_EN_clint_mtime = EN_clint_mtime ;
  assign csr_EN_incr_minstret = WILL_FIRE_RL_increment_instruction_counter ;
  assign csr_EN_ext_interrupt = EN_ext_interrupt ;

  // submodule dump_ff
  assign dump_ff_D_IN =
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179) ?
	       { IF_csr_mv_curr_priv__83_EQ_3_84_THEN_csr_mv_cu_ETC___d185,
		 rx_stage3_dump_first_x,
		 rx_stage3_common_first_x[5:1],
		 data__h3311 } :
	       _dfoo2 ;
  assign dump_ff_ENQ =
	     WILL_FIRE_RL_instruction_commit &&
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 ||
	      _dfoo1) ;
  assign dump_ff_DEQ = EN_dump_get ;
  assign dump_ff_CLR = 1'b0 ;

  // remaining internal signals
  assign IF_csr_mv_curr_priv__83_EQ_3_84_THEN_csr_mv_cu_ETC___d185 =
	     (csr_mv_curr_priv == 2'd3) ? csr_mv_curr_priv : 2'd0 ;
  assign IF_ff_stage3_dump_w_data_whas__5_THEN_ff_stage_ETC___d237 =
	     { rx_stage3_dump_first_x[31:0],
	       (IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
		2'd2) ?
		 69'd0 :
		 { rx_stage3_common_first_x[5:1], _theResult____h4431 } } ;
  assign NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 =
	     !rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd2 &&
	     (!ff_stage3_type_w_data_wget[0] || ma_delayed_output_r[0]) ;
  assign NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190 =
	     !rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd2 &&
	     ff_stage3_type_w_data_wget[0] &&
	     !ma_delayed_output_r[0] ;
  assign NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202 =
	     !rg_rerun && ff_stage3_type_w_data_wget[82:81] != 2'd0 &&
	     ff_stage3_type_w_data_wget[82:81] != 2'd1 &&
	     ff_stage3_type_w_data_wget[82:81] != 2'd2 ;
  assign _dfoo1 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     (NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202 ||
	      !rg_rerun &&
	      ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d224) ;
  assign _dfoo10 =
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202) ?
	       { 1'd1, rx_stage3_common_first_x[5:1], _theResult____h4120 } :
	       ((IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
		 2'd2) ?
		  70'h200000000000000000 :
		  { 1'd1,
		    rx_stage3_common_first_x[5:1],
		    _theResult____h4431 }) ;
  assign _dfoo14 =
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      !rg_rerun &&
	      ff_stage3_type_w_data_whas__1_AND_NOT_ff_stage_ETC___d204) ?
	       { csr_system_instruction[127:64], 1'd1 } :
	       { csr_take_trap, 1'd1 } ;
  assign _dfoo2 =
	     (rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	      NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202) ?
	       { IF_csr_mv_curr_priv__83_EQ_3_84_THEN_csr_mv_cu_ETC___d185,
		 rx_stage3_dump_first_x,
		 rx_stage3_common_first_x[5:1],
		 _theResult____h4120 } :
	       { IF_csr_mv_curr_priv__83_EQ_3_84_THEN_csr_mv_cu_ETC___d185,
		 rx_stage3_dump_first_x[95:32],
		 IF_ff_stage3_dump_w_data_whas__5_THEN_ff_stage_ETC___d237 } ;
  assign _dfoo25 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d164 ||
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     !rg_rerun &&
	     ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	     IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 !=
	     2'd2 &&
	     wr_memory_response[66] &&
	     wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218 &&
	     !wr_memory_response[1] ;
  assign _dfoo3 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     (NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d202 ||
	      !rg_rerun &&
	      ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d233) ;
  assign _dfoo31 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     (rg_rerun ||
	      ff_stage3_type_w_data_wget[82:81] != 2'd0 &&
	      ff_stage3_type_w_data_wget[82:81] != 2'd1 &&
	      ff_stage3_type_w_data_wget[82:81] != 2'd2 &&
	      !csr_system_instruction[128] ||
	      !rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	      IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
	      2'd2) ;
  assign _dfoo33 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d128 ||
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     !rg_rerun &&
	     (ff_stage3_type_w_data_whas__1_AND_NOT_ff_stage_ETC___d204 ||
	      ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243) ;
  assign _dfoo37 =
	     rg_rerun_22_OR_ff_stage3_type_w_data_whas__1_A_ETC___d127 ||
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 ||
	     _dfoo3 ;
  assign _dfoo39 =
	     rg_rerun_22_OR_ff_stage3_type_w_data_whas__1_A_ETC___d127 ||
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 ||
	     _dfoo3 ;
  assign _dfoo41 =
	     rg_rerun_22_OR_ff_stage3_type_w_data_whas__1_A_ETC___d127 ||
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d179 ||
	     _dfoo3 ;
  assign _theResult_____1_snd__h3364 =
	     (!ma_delayed_output_r[0] ||
	      rx_stage3_common_first_x[5:1] == 5'd0) ?
	       _theResult____h3307 :
	       ma_delayed_output_r[64:1] ;
  assign _theResult____h3307 =
	     (rx_stage3_common_first_x[5:1] == 5'd0) ?
	       64'd0 :
	       ff_stage3_type_w_data_wget[64:1] ;
  assign _theResult____h4120 =
	     (rx_stage3_common_first_x[5:1] == 5'd0) ?
	       64'd0 :
	       csr_system_instruction[63:0] ;
  assign _theResult____h4431 =
	     (rx_stage3_common_first_x[5:1] == 5'd0) ?
	       64'd0 :
	       wr_memory_response[65:2] ;
  assign data__h3311 =
	     ff_stage3_type_w_data_wget[0] ?
	       _theResult_____1_snd__h3364 :
	       _theResult____h3307 ;
  assign ff_stage3_type_w_data_whas__1_AND_NOT_ff_stage_ETC___d204 =
	     ff_stage3_type_w_data_wget[82:81] != 2'd0 &&
	     ff_stage3_type_w_data_wget[82:81] != 2'd1 &&
	     ff_stage3_type_w_data_wget[82:81] != 2'd2 &&
	     csr_system_instruction[128] ;
  assign ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d224 =
	     ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	     (IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
	      2'd2 ||
	      wr_memory_response[66] &&
	      wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218 &&
	      !wr_memory_response[1]) ;
  assign ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d233 =
	     ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	     (IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
	      2'd2 ||
	      wr_memory_response[66] &&
	      wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218) ;
  assign ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243 =
	     ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	     IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 !=
	     2'd2 &&
	     wr_memory_response[66] &&
	     wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218 &&
	     wr_memory_response[1] ;
  assign ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269 =
	     ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	     IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 !=
	     2'd2 &&
	     (!wr_memory_response[66] ||
	      !wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218) ;
  assign rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 =
	     rg_epoch == rx_stage3_common_first_x[0] ;
  assign rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d128 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     (rg_rerun || ff_stage3_type_w_data_wget[82:81] == 2'd1) ;
  assign rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     !rg_rerun &&
	     ff_stage3_type_w_data_wget[82:81] == 2'd1 ;
  assign rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d164 =
	     rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	     !rg_rerun &&
	     ff_stage3_type_w_data_wget[82:81] == 2'd2 ;
  assign rg_rerun_22_OR_ff_stage3_type_w_data_whas__1_A_ETC___d127 =
	     rg_rerun || ff_stage3_type_w_data_wget[82:81] == 2'd1 ||
	     !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 ;
  assign type_cause__h4513 =
	     (IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 ==
	      2'd0) ?
	       6'd5 :
	       6'd7 ;
  assign wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218 =
	     wr_memory_response[0] == rg_epoch ;
  assign x__h4837 = ~rg_epoch ;
  assign x__read_rdaddr__h5758 =
	     wr_operand_fwding_whas ? wr_operand_fwding_wget[69:65] : 5'd0 ;
  assign x__read_rdvalue__h5759 =
	     wr_operand_fwding_whas ? wr_operand_fwding_wget[64:1] : 64'd0 ;
  always@(csr_mv_trigger_data1)
  begin
    case (csr_mv_trigger_data1[43:42])
      2'd0, 2'd1, 2'd2:
	  CASE_csrmv_trigger_data1_BITS_43_TO_42_0_csr_ETC__q1 =
	      csr_mv_trigger_data1[43:22];
      2'd3:
	  CASE_csrmv_trigger_data1_BITS_43_TO_42_0_csr_ETC__q1 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(csr_mv_trigger_data1)
  begin
    case (csr_mv_trigger_data1[21:20])
      2'd0, 2'd1, 2'd2:
	  CASE_csrmv_trigger_data1_BITS_21_TO_20_0_csr_ETC__q2 =
	      csr_mv_trigger_data1[21:0];
      2'd3:
	  CASE_csrmv_trigger_data1_BITS_21_TO_20_0_csr_ETC__q2 =
	      { 2'd3, 20'b10101010101010101010 /* unspecified value */  };
    endcase
  end
  always@(rx_stage3_type_first_x)
  begin
    case (rx_stage3_type_first_x[82:81])
      2'd0, 2'd1, 2'd2:
	  CASE_rx_stage3_type_first_x_BITS_82_TO_81_0_rx_ETC__q3 =
	      rx_stage3_type_first_x[82:81];
      2'd3: CASE_rx_stage3_type_first_x_BITS_82_TO_81_0_rx_ETC__q3 = 2'd3;
    endcase
  end
  always@(rx_stage3_type_first_x)
  begin
    case (rx_stage3_type_first_x[67:66])
      2'd0, 2'd1, 2'd3:
	  CASE_rx_stage3_type_first_x_BITS_67_TO_66_0_rx_ETC__q4 =
	      rx_stage3_type_first_x[67:66];
      2'd2: CASE_rx_stage3_type_first_x_BITS_67_TO_66_0_rx_ETC__q4 = 2'd2;
    endcase
  end
  always@(ff_stage3_type_w_data_wget)
  begin
    case (ff_stage3_type_w_data_wget[67:66])
      2'd0, 2'd1:
	  IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 =
	      ff_stage3_type_w_data_wget[67:66];
      2'd2: IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 = 2'd3;
      2'd3: IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 = 2'd2;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_epoch <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_rerun <= `BSV_ASSIGNMENT_DELAY 1'd0;
	wr_memory_response <= `BSV_ASSIGNMENT_DELAY
	    { 1'd0, 66'h2AAAAAAAAAAAAAAAA /* unspecified value */  };
      end
    else
      begin
        if (rg_epoch_EN) rg_epoch <= `BSV_ASSIGNMENT_DELAY rg_epoch_D_IN;
	if (rg_rerun_EN) rg_rerun <= `BSV_ASSIGNMENT_DELAY rg_rerun_D_IN;
	if (wr_memory_response_EN)
	  wr_memory_response <= `BSV_ASSIGNMENT_DELAY wr_memory_response_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_epoch = 1'h0;
    rg_rerun = 1'h0;
    wr_memory_response = 67'h2AAAAAAAAAAAAAAAA;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d19 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d20 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d21 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  v__h1870 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("[%10d", v__h1870, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("STAGE3: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("TraceDump { ", "pc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("'h%h", rx_stage3_dump_first_x[95:32]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write(", ", "instruction: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("'h%h", rx_stage3_dump_first_x[31:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d19 ||
	   TASK_testplusargs___d20 && TASK_testplusargs___d21))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d31 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d32 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d33 = $test$plusargs("l0");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  v__h2055 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("[%10d", v__h2055, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("STAGE3: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("Stage3Common { ", "pc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("'h%h", rx_stage3_common_first_x[69:6]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write(", ", "rd: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("'h%h", rx_stage3_common_first_x[5:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write(", ", "epoch: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("'h%h", rx_stage3_common_first_x[0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d31 ||
	   TASK_testplusargs___d32 && TASK_testplusargs___d33))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d45 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d46 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  TASK_testplusargs___d47 = $test$plusargs("l0");
	  #0;
	end
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd0;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd1;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd2;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] != 2'd0 &&
	ff_stage3_type_w_data_wget[82:81] != 2'd1 &&
	ff_stage3_type_w_data_wget[82:81] != 2'd2;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d85 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd2 &&
	ff_stage3_type_w_data_wget[0];
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d88 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd2 &&
	!ff_stage3_type_w_data_wget[0];
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] != 2'd0 &&
	ff_stage3_type_w_data_wget[82:81] != 2'd1;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] != 2'd0;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d106 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 == 2'd0;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d109 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 == 2'd1;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d112 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 == 2'd2;
    TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d119 =
	(TASK_testplusargs___d45 ||
	 TASK_testplusargs___d46 && TASK_testplusargs___d47) &&
	ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 != 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 != 2'd1 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 != 2'd2;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit)
	begin
	  v__h2250 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d45 ||
	   TASK_testplusargs___d46 && TASK_testplusargs___d47))
	$write("[%10d", v__h2250, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d45 ||
	   TASK_testplusargs___d46 && TASK_testplusargs___d47))
	$write("STAGE3: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("tagged Memory ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("tagged Trap ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("tagged Regular ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("tagged System ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("Stage3System { ", "rs1_imm: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("'h%h", ff_stage3_type_w_data_wget[80:17]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write(", ", "lpc: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("'h%h", ff_stage3_type_w_data_wget[16:15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write(", ", "csr_address: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("'h%h", ff_stage3_type_w_data_wget[14:3]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write(", ", "funct3: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("'h%h", ff_stage3_type_w_data_wget[2:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("Stage3Regular { ", "rdvalue: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write("'h%h", ff_stage3_type_w_data_wget[64:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write(", ", "delayed: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d85)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d88)
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d62)
	$write(" }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d72)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("Stage3Trap { ", "cause: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("'h%h", ff_stage3_type_w_data_wget[69:64]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write(", ", "badaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d59)
	$write("'h%h", ff_stage3_type_w_data_wget[63:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d90)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("Stage3Memory { ", "memaccess: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d106)
	$write("Load");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d109)
	$write("Store");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d112)
	$write("Fence");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d119)
	$write("Atomic");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write(", ", "address: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("'h%h", ff_stage3_type_w_data_wget[65:2]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write(", ", "size: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d56)
	$write("'h%h", ff_stage3_type_w_data_wget[1:0], " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  TASK_testplusargs_5_OR_TASK_testplusargs_6_AND_ETC___d95)
	$write("");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  (TASK_testplusargs___d45 ||
	   TASK_testplusargs___d46 && TASK_testplusargs___d47))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun)
	begin
	  TASK_testplusargs___d144 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun)
	begin
	  TASK_testplusargs___d145 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun)
	begin
	  TASK_testplusargs___d146 = $test$plusargs("l0");
	  #0;
	end
    rg_rerun_22_AND_TASK_testplusargs_44_OR_TASK_t_ETC___d149 =
	rg_rerun &&
	(TASK_testplusargs___d144 ||
	 TASK_testplusargs___d145 && TASK_testplusargs___d146);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun)
	begin
	  v__h3248 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun_22_AND_TASK_testplusargs_44_OR_TASK_t_ETC___d149)
	$write("[%10d", v__h3248, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun_22_AND_TASK_testplusargs_44_OR_TASK_t_ETC___d149)
	$write("STAGE3: Rerun Instruction");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  rg_rerun_22_AND_TASK_testplusargs_44_OR_TASK_t_ETC___d149)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153)
	begin
	  TASK_testplusargs___d154 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153)
	begin
	  TASK_testplusargs___d155 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153)
	begin
	  TASK_testplusargs___d156 = $test$plusargs("l0");
	  #0;
	end
    ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d159 =
	ff_stage3_type_w_data_wget[82:81] == 2'd1 &&
	(TASK_testplusargs___d154 ||
	 TASK_testplusargs___d155 && TASK_testplusargs___d156);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d153)
	begin
	  v__h2907 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d159)
	$write("[%10d", v__h2907, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d159)
	$write("STAGE3 : Jumping to PC:%h", csr_take_trap);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d159)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190)
	begin
	  TASK_testplusargs___d192 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190)
	begin
	  TASK_testplusargs___d193 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190)
	begin
	  TASK_testplusargs___d194 = $test$plusargs("l0");
	  #0;
	end
    ff_stage3_type_w_data_wget__2_BIT_0_3_AND_NOT__ETC___d197 =
	ff_stage3_type_w_data_wget[0] && !ma_delayed_output_r[0] &&
	(TASK_testplusargs___d192 ||
	 TASK_testplusargs___d193 && TASK_testplusargs___d194);
    NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d199 =
	!rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd2 &&
	ff_stage3_type_w_data_wget__2_BIT_0_3_AND_NOT__ETC___d197;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d190)
	begin
	  v__h3730 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d199)
	$write("[%10d", v__h3730, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d199)
	$write("STAGE3: Waiting for Delayed Output");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d199)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243)
	begin
	  TASK_testplusargs___d248 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243)
	begin
	  TASK_testplusargs___d249 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243)
	begin
	  TASK_testplusargs___d250 = $test$plusargs("l0");
	  #0;
	end
    wr_memory_response_15_BIT_1_20_AND_TASK_testpl_ETC___d253 =
	wr_memory_response[1] &&
	(TASK_testplusargs___d248 ||
	 TASK_testplusargs___d249 && TASK_testplusargs___d250);
    NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d257 =
	!rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 != 2'd2 &&
	wr_memory_response[66] &&
	wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218 &&
	wr_memory_response_15_BIT_1_20_AND_TASK_testpl_ETC___d253;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d243)
	begin
	  v__h4969 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d257)
	$write("[%10d", v__h4969, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d257)
	$write("STAGE3 : Jumping to PC:%h", csr_take_trap);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d257)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269)
	begin
	  TASK_testplusargs___d272 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269)
	begin
	  TASK_testplusargs___d273 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269)
	begin
	  TASK_testplusargs___d274 = $test$plusargs("l1");
	  #0;
	end
    NOT_wr_memory_response_15_BIT_66_16_65_OR_NOT__ETC___d277 =
	(!wr_memory_response[66] ||
	 !wr_memory_response_15_BIT_0_17_EQ_rg_epoch_24___d218) &&
	(TASK_testplusargs___d272 ||
	 TASK_testplusargs___d273 && TASK_testplusargs___d274);
    NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d280 =
	!rg_rerun && ff_stage3_type_w_data_wget[82:81] == 2'd0 &&
	IF_ff_stage3_type_w_data_whas__1_THEN_IF_ff_st_ETC___d103 != 2'd2 &&
	NOT_wr_memory_response_15_BIT_66_16_65_OR_NOT__ETC___d277;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  !rg_rerun &&
	  ff_stage3_type_w_data_whas__1_AND_ff_stage3_ty_ETC___d269)
	begin
	  v__h5043 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d280)
	$write("[%10d", v__h5043, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d280)
	$write("STAGE3 : Waiting for response from Fabric");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	  NOT_rg_rerun_22_42_AND_ff_stage3_type_w_data_w_ETC___d280)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125)
	begin
	  TASK_testplusargs___d283 = $test$plusargs("fullverbose");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125)
	begin
	  TASK_testplusargs___d284 = $test$plusargs("mstage3");
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125)
	begin
	  TASK_testplusargs___d285 = $test$plusargs("l0");
	  #0;
	end
    NOT_rg_epoch_24_EQ_IF_ff_stage3_common_w_data__ETC___d288 =
	!rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125 &&
	(TASK_testplusargs___d283 ||
	 TASK_testplusargs___d284 && TASK_testplusargs___d285);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  !rg_epoch_24_EQ_IF_ff_stage3_common_w_data_whas_ETC___d125)
	begin
	  v__h5138 = $time;
	  #0;
	end
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  NOT_rg_epoch_24_EQ_IF_ff_stage3_common_w_data__ETC___d288)
	$write("[%10d", v__h5138, "] ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  NOT_rg_epoch_24_EQ_IF_ff_stage3_common_w_data__ETC___d288)
	$write("STAGE3 : Dropping instruction");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_instruction_commit &&
	  NOT_rg_epoch_24_EQ_IF_ff_stage3_common_w_data__ETC___d288)
	$write("\n");
  end
  // synopsys translate_on
endmodule  // mkstage3

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:51 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// CLK                            I     1 unused
// RST_N                          I     1 unused
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkTb(CLK,
	    RST_N);
  input  CLK;
  input  RST_N;

endmodule  // mkTb

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:53 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// address_valid                  O     1
// address_valid_addr             I    12
// address_valid_misa             I    26
//
// Combinational paths from inputs to outputs:
//   (address_valid_addr, address_valid_misa) -> address_valid
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_address_valid(address_valid_addr,
			    address_valid_misa,
			    address_valid);
  // value method address_valid
  input  [11 : 0] address_valid_addr;
  input  [25 : 0] address_valid_misa;
  output address_valid;

  // signals for module outputs
  wire address_valid;

  // remaining internal signals
  reg CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q2,
      CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5,
      CASE_address_valid_addr_BITS_7_TO_0_0_address__ETC__q1,
      CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4,
      CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3;
  wire address_valid_addr_BITS_3_TO_0_0_EQ_0x0_0_OR_a_ETC___d61,
       address_valid_misa_BIT_13_1_AND_address_valid__ETC___d23;

  // value method address_valid
  assign address_valid =
	     (address_valid_addr[9:8] == 2'b0) ?
	       CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q2 :
	       address_valid_addr[9:8] == 2'b11 &&
	       CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5 ;

  // remaining internal signals
  assign address_valid_addr_BITS_3_TO_0_0_EQ_0x0_0_OR_a_ETC___d61 =
	     address_valid_addr[3:0] == 4'h0 ||
	     address_valid_addr[3:0] == 4'd1 ||
	     address_valid_addr[3:0] == 4'h4 ||
	     address_valid_addr[3:0] == 4'h5 ||
	     address_valid_addr[3:0] == 4'h6 ||
	     (address_valid_addr[3:0] == 4'h2 ||
	      address_valid_addr[3:0] == 4'h3) &&
	     (address_valid_misa_BIT_13_1_AND_address_valid__ETC___d23 ||
	      address_valid_misa[18]) ;
  assign address_valid_misa_BIT_13_1_AND_address_valid__ETC___d23 =
	     address_valid_misa[13] & address_valid_misa[20] ;
  always@(address_valid_addr or
	  address_valid_misa_BIT_13_1_AND_address_valid__ETC___d23)
  begin
    case (address_valid_addr[7:0])
      8'd0, 8'h04, 8'h05, 8'h40, 8'h41, 8'h42, 8'h43, 8'h44:
	  CASE_address_valid_addr_BITS_7_TO_0_0_address__ETC__q1 =
	      address_valid_misa_BIT_13_1_AND_address_valid__ETC___d23;
      default: CASE_address_valid_addr_BITS_7_TO_0_0_address__ETC__q1 =
		   address_valid_addr[7:0] == 8'h01 ||
		   address_valid_addr[7:0] == 8'h02 ||
		   address_valid_addr[7:0] == 8'h03;
    endcase
  end
  always@(address_valid_addr or
	  CASE_address_valid_addr_BITS_7_TO_0_0_address__ETC__q1)
  begin
    case (address_valid_addr[11:10])
      2'b0:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q2 =
	      CASE_address_valid_addr_BITS_7_TO_0_0_address__ETC__q1;
      2'b11:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q2 =
	      address_valid_addr[7:5] == 3'b0;
      default: CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q2 =
		   address_valid_addr[11:10] == 2'b10 &&
		   address_valid_addr[7:0] == 8'd0;
    endcase
  end
  always@(address_valid_addr)
  begin
    case (address_valid_addr[7:4])
      4'h4:
	  CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3 =
	      address_valid_addr[3:0] == 4'h0 ||
	      address_valid_addr[3:0] == 4'd1 ||
	      address_valid_addr[3:0] == 4'h2 ||
	      address_valid_addr[3:0] == 4'h3 ||
	      address_valid_addr[3:0] == 4'h4;
      4'hA:
	  CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3 =
	      address_valid_addr[3:0] == 4'h0 ||
	      address_valid_addr[3:0] == 4'h2;
      default: CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3 =
		   address_valid_addr[7:4] == 4'hB &&
		   address_valid_addr[3:0] <= 4'd3;
    endcase
  end
  always@(address_valid_addr or
	  CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3 or
	  address_valid_addr_BITS_3_TO_0_0_EQ_0x0_0_OR_a_ETC___d61)
  begin
    case (address_valid_addr[7:4])
      4'd0:
	  CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4 =
	      address_valid_addr_BITS_3_TO_0_0_EQ_0x0_0_OR_a_ETC___d61;
      4'h2:
	  CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4 =
	      address_valid_addr[3:0] > 4'd2;
      default: CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4 =
		   address_valid_addr[7:4] == 4'h3 ||
		   CASE_address_valid_addr_BITS_7_TO_4_0x4_addres_ETC__q3;
    endcase
  end
  always@(address_valid_addr or
	  CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4)
  begin
    case (address_valid_addr[11:10])
      2'b0:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5 =
	      CASE_address_valid_addr_BITS_7_TO_4_0_address__ETC__q4;
      2'd1:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5 =
	      address_valid_addr[11:10] == 2'b01 &&
	      address_valid_addr[7:4] == 4'hA &&
	      address_valid_addr[3:0] < 4'd4;
      2'b10:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5 =
	      address_valid_addr[7:4] == 4'd0 &&
	      address_valid_addr[3:0] != 4'd1;
      2'b11:
	  CASE_address_valid_addr_BITS_11_TO_10_0b0_CASE_ETC__q5 =
	      address_valid_addr[7:4] == 4'd1 &&
	      (address_valid_addr[3:0] == 4'd1 ||
	       address_valid_addr[3:0] == 4'h2 ||
	       address_valid_addr[3:0] == 4'h3 ||
	       address_valid_addr[3:0] == 4'h4);
    endcase
  end
endmodule  // module_address_valid

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:53 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// chk_interrupt                  O     8
// chk_interrupt_prv              I     2
// chk_interrupt_mstatus          I    64
// chk_interrupt_mip              I    14
// chk_interrupt_mie              I    12
// chk_interrupt_mideleg          I    12
// chk_interrupt_uip              I    12
// chk_interrupt_uie              I    12
//
// Combinational paths from inputs to outputs:
//   (chk_interrupt_prv,
//    chk_interrupt_mstatus,
//    chk_interrupt_mip,
//    chk_interrupt_mie,
//    chk_interrupt_mideleg,
//    chk_interrupt_uip,
//    chk_interrupt_uie) -> chk_interrupt
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_chk_interrupt(chk_interrupt_prv,
			    chk_interrupt_mstatus,
			    chk_interrupt_mip,
			    chk_interrupt_mie,
			    chk_interrupt_mideleg,
			    chk_interrupt_uip,
			    chk_interrupt_uie,
			    chk_interrupt);
  // value method chk_interrupt
  input  [1 : 0] chk_interrupt_prv;
  input  [63 : 0] chk_interrupt_mstatus;
  input  [13 : 0] chk_interrupt_mip;
  input  [11 : 0] chk_interrupt_mie;
  input  [11 : 0] chk_interrupt_mideleg;
  input  [11 : 0] chk_interrupt_uip;
  input  [11 : 0] chk_interrupt_uie;
  output [7 : 0] chk_interrupt;

  // signals for module outputs
  wire [7 : 0] chk_interrupt;

  // remaining internal signals
  wire [13 : 0] pending_interrupts__h39;
  wire [11 : 0] m_interrupts__h37,
		u_interrupts__h38,
		x__h155,
		x__h209,
		x__h211,
		x__h350,
		y__h156,
		y__h158,
		y__h210;
  wire [5 : 0] x__h28;

  // value method chk_interrupt
  assign chk_interrupt =
	     { x__h28, pending_interrupts__h39 != 14'd0, x__h350 != 12'd0 } ;

  // remaining internal signals
  assign m_interrupts__h37 = x__h155 & y__h156 ;
  assign pending_interrupts__h39 =
	     ((chk_interrupt_prv != 2'd3 || chk_interrupt_mstatus[3]) ?
		{ 2'd0, m_interrupts__h37 } :
		14'd0) |
	     ((chk_interrupt_mstatus[0] && chk_interrupt_prv != 2'd3) ?
		{ 2'd0, u_interrupts__h38 } :
		14'd0) ;
  assign u_interrupts__h38 = x__h209 & y__h210 ;
  assign x__h155 = x__h350 & y__h158 ;
  assign x__h209 = x__h211 & chk_interrupt_mideleg ;
  assign x__h211 = chk_interrupt_uie & chk_interrupt_uip ;
  assign x__h28 =
	     { 1'b1,
	       pending_interrupts__h39[11] ?
		 5'd11 :
		 (pending_interrupts__h39[3] ?
		    5'd3 :
		    (pending_interrupts__h39[7] ?
		       5'd7 :
		       (pending_interrupts__h39[8] ?
			  5'd8 :
			  (pending_interrupts__h39[0] ?
			     5'd0 :
			     (pending_interrupts__h39[4] ?
				5'd4 :
				5'd31))))) } ;
  assign x__h350 = chk_interrupt_mie & chk_interrupt_mip[11:0] ;
  assign y__h156 = ~chk_interrupt_mideleg ;
  assign y__h158 =
	     {12{chk_interrupt_prv != 2'd3 || chk_interrupt_mstatus[3]}} ;
  assign y__h210 =
	     {12{chk_interrupt_mstatus[0] && chk_interrupt_prv != 2'd3}} ;
endmodule  // module_chk_interrupt

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:53 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// decoder_func_32                O    65
// decoder_func_32_inst           I    32
// decoder_func_32_csrs           I   152
// decoder_func_32_compressed     I     1
//
// Combinational paths from inputs to outputs:
//   (decoder_func_32_inst,
//    decoder_func_32_csrs,
//    decoder_func_32_compressed) -> decoder_func_32
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_decoder_func_32(decoder_func_32_inst,
			      decoder_func_32_csrs,
			      decoder_func_32_compressed,
			      decoder_func_32);
  // value method decoder_func_32
  input  [31 : 0] decoder_func_32_inst;
  input  [151 : 0] decoder_func_32_csrs;
  input  decoder_func_32_compressed;
  output [64 : 0] decoder_func_32;

  // signals for module outputs
  wire [64 : 0] decoder_func_32;

  // remaining internal signals
  reg [10 : 0] CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q10;
  reg [7 : 0] CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q11;
  reg [5 : 0] CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q8,
	      _theResult_____6_snd__h1554,
	      _theResult_____6_snd__h1609;
  reg [4 : 0] x__h268;
  reg [3 : 0] CASE_decoder_func_32_inst_BITS_14_TO_12_0_1_1_1_6__q12,
	      CASE_decoder_func_32_inst_BITS_31_TO_7_0_6_0x2_ETC__q1,
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14,
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13,
	      CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q9,
	      CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15,
	      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212,
	      IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432,
	      fn___1__h4966,
	      fn___1__h5028;
  reg [1 : 0] CASE_decoder_func_32_inst_BITS_6_TO_2_0b0_1_0b_ETC__q17,
	      CASE_decoder_func_32_inst_BITS_6_TO_2_0b11_3_0_ETC__q16;
  reg CASE_decoder_func_32_inst_BITS_14_TO_12_0_NOT__ETC__q5,
      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2,
      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3,
      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6,
      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7,
      CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q4,
      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119,
      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132,
      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301,
      IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337;
  wire [41 : 0] IF_NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1_ETC___d436;
  wire [31 : 0] immediate_value___1__h2154,
		immediate_value__h49,
		instr_meta_immediate__h351;
  wire [11 : 0] NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1011_ETC___d371;
  wire [10 : 0] bit20_30__h47;
  wire [7 : 0] bit12_19__h46;
  wire [6 : 0] instr_meta_funct__h352, temp1___1__h4863, temp1__h70;
  wire [5 : 0] _theResult_____6_snd__h1582, trapcause___1__h1604, x__h4866;
  wire [4 : 0] x__h194, x__h21;
  wire [3 : 0] IF_NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0_ETC___d228,
	       IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d205,
	       IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d207,
	       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d220,
	       IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411,
	       fn___1__h4927,
	       fn___1__h4949;
  wire [1 : 0] IF_decoder_func_32_compressed_THEN_3_ELSE_2___d40;
  wire IF_decoder_func_32_csrs_BITS_151_TO_150_55_EQ__ETC___d169,
       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d184,
       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d330,
       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d340,
       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d126,
       IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68,
       NOT_decoder_func_32_csrs_BIT_76_15_86_OR_NOT_d_ETC___d296,
       NOT_decoder_func_32_inst_BITS_14_TO_12_3_EQ_4__ETC___d180,
       NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0b11_ETC___d192,
       address_valid___d182,
       bit31__h48,
       decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114,
       decoder_func_32_csrs_BIT_76_15_AND_decoder_fun_ETC___d127,
       decoder_func_32_inst_BITS_14_TO_12_3_ULE_3___d121,
       decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84,
       decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158,
       decoder_func_32_inst_BIT_27_21_OR_decoder_func_ETC___d423;

  // value method decoder_func_32
  assign decoder_func_32 =
	     { x__h21,
	       x__h194,
	       x__h268,
	       decoder_func_32_inst[6:2] == 5'b11011 ||
	       decoder_func_32_inst[6:2] == 5'b11001 ||
	       decoder_func_32_inst[6:2] == 5'b00101,
	       CASE_decoder_func_32_inst_BITS_6_TO_2_0b0_1_0b_ETC__q17,
	       IF_NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0_ETC___d228,
	       IF_NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1_ETC___d436,
	       1'd0 } ;

  // remaining internal signals
  module_address_valid instance_address_valid_0(.address_valid_addr(decoder_func_32_inst[31:20]),
						.address_valid_misa(decoder_func_32_csrs[89:64]),
						.address_valid(address_valid___d182));
  assign IF_NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0_ETC___d228 =
	     NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0b11_ETC___d192 ?
	       4'd6 :
	       CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15 ;
  assign IF_NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1_ETC___d436 =
	     { (decoder_func_32_inst[6:2] != 5'b01011 &&
		decoder_func_32_inst[6:2] != 5'b00011 &&
		decoder_func_32_inst[6:2] != 5'b01000) ?
		 2'd0 :
		 CASE_decoder_func_32_inst_BITS_6_TO_2_0b11_3_0_ETC__q16,
	       instr_meta_immediate__h351,
	       instr_meta_funct__h352,
	       1'b0 /* unspecified value */  } ;
  assign IF_decoder_func_32_compressed_THEN_3_ELSE_2___d40 =
	     decoder_func_32_compressed ? 2'd3 : 2'd2 ;
  assign IF_decoder_func_32_csrs_BITS_151_TO_150_55_EQ__ETC___d169 =
	     ((decoder_func_32_csrs[151:150] == 2'd3) ?
		decoder_func_32_csrs[151:150] :
		2'd0) <
	     decoder_func_32_inst[29:28] ;
  assign IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d205 =
	     (decoder_func_32_csrs[76] &&
	      decoder_func_32_inst[31:25] == 7'd1) ?
	       4'd8 :
	       (IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119 ?
		  4'd0 :
		  4'd6) ;
  assign IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d207 =
	     (decoder_func_32_csrs[76] &&
	      decoder_func_32_inst[31:25] == 7'd1 &&
	      (decoder_func_32_inst[14:12] == 3'd0 ||
	       !decoder_func_32_inst_BITS_14_TO_12_3_ULE_3___d121)) ?
	       4'd8 :
	       (IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d126 ?
		  4'd0 :
		  4'd6) ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d184 =
	     (decoder_func_32_inst[14:12] == 3'd0) ?
	       decoder_func_32_inst[31:7] != 25'd0 &&
	       decoder_func_32_inst[31:7] != 25'h0002000 &&
	       (decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158 ||
		decoder_func_32_inst[31:20] == 12'h105 &&
		decoder_func_32_inst[19:15] == 5'd0 &&
		decoder_func_32_inst[11:7] == 5'd0 &&
		decoder_func_32_csrs[151:150] == 2'd3) :
	       NOT_decoder_func_32_inst_BITS_14_TO_12_3_EQ_4__ETC___d180 &&
	       address_valid___d182 ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d220 =
	     (decoder_func_32_inst[14:12] == 3'd0) ?
	       CASE_decoder_func_32_inst_BITS_31_TO_7_0_6_0x2_ETC__q1 :
	       ((NOT_decoder_func_32_inst_BITS_14_TO_12_3_EQ_4__ETC___d180 &&
		 address_valid___d182) ?
		  4'd5 :
		  4'd6) ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d330 =
	     (decoder_func_32_inst[14:12] == 3'd0) ?
	       (decoder_func_32_inst[31:20] != 12'h002 ||
		decoder_func_32_inst[19:15] != 5'd0 ||
		decoder_func_32_inst[11:7] != 5'd0 ||
		!decoder_func_32_csrs[77]) &&
	       (decoder_func_32_inst[31:20] != 12'h302 ||
		decoder_func_32_inst[19:15] != 5'd0 ||
		decoder_func_32_inst[11:7] != 5'd0 ||
		decoder_func_32_csrs[151:150] != 2'd3) &&
	       (decoder_func_32_inst[31:20] != 12'h105 ||
		decoder_func_32_inst[19:15] != 5'd0 ||
		decoder_func_32_inst[11:7] != 5'd0 ||
		decoder_func_32_csrs[151:150] != 2'd3) :
	       decoder_func_32_inst[14:12] == 3'd4 ||
	       IF_decoder_func_32_csrs_BITS_151_TO_150_55_EQ__ETC___d169 ||
	       (decoder_func_32_inst[19:15] != 5'd0 ||
		decoder_func_32_inst[13:12] == 2'b01) &&
	       decoder_func_32_inst[31:30] == 2'b11 ||
	       !address_valid___d182 ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d340 =
	     (decoder_func_32_inst[14:12] == 3'd0) ?
	       decoder_func_32_inst[31:7] != 25'd0 &&
	       decoder_func_32_inst[31:7] != 25'h0002000 &&
	       decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158 :
	       NOT_decoder_func_32_inst_BITS_14_TO_12_3_EQ_4__ETC___d180 &&
	       address_valid___d182 ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d126 =
	     (decoder_func_32_inst[14:12] == 3'd1) ?
	       decoder_func_32_inst[31:25] == 7'b0 :
	       (decoder_func_32_inst[14:12] == 3'd0 ||
		decoder_func_32_inst[14:12] == 3'd5) &&
	       (decoder_func_32_inst[31:25] == 7'b0 ||
		decoder_func_32_inst[31:25] == 7'b0100000) ;
  assign IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68 =
	     (decoder_func_32_inst[14:12] == 3'd1) ?
	       decoder_func_32_inst[31:26] == 6'd0 :
	       decoder_func_32_inst[14:12] != 3'd5 ||
	       decoder_func_32_inst[31:26] == 6'd0 ||
	       decoder_func_32_inst[31:26] == 6'b010000 ;
  assign IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411 =
	     decoder_func_32_inst[30] ? 4'b1011 : 4'b0101 ;
  assign NOT_decoder_func_32_csrs_BIT_76_15_86_OR_NOT_d_ETC___d296 =
	     (!decoder_func_32_csrs[76] ||
	      decoder_func_32_inst[31:25] != 7'd1 ||
	      decoder_func_32_inst[14:12] != 3'd0 &&
	      decoder_func_32_inst_BITS_14_TO_12_3_ULE_3___d121) &&
	     ((decoder_func_32_inst[14:12] == 3'd1) ?
		decoder_func_32_inst[31:25] != 7'b0 :
		decoder_func_32_inst[14:12] != 3'd0 &&
		decoder_func_32_inst[14:12] != 3'd5 ||
		decoder_func_32_inst[31:25] != 7'b0 &&
		decoder_func_32_inst[31:25] != 7'b0100000) ;
  assign NOT_decoder_func_32_inst_BITS_14_TO_12_3_EQ_4__ETC___d180 =
	     decoder_func_32_inst[14:12] != 3'd4 &&
	     !IF_decoder_func_32_csrs_BITS_151_TO_150_55_EQ__ETC___d169 &&
	     (decoder_func_32_inst[19:15] == 5'd0 &&
	      decoder_func_32_inst[13:12] != 2'b01 ||
	      decoder_func_32_inst[31:30] != 2'b11) ;
  assign NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0b11_ETC___d192 =
	     decoder_func_32_inst[1:0] != 2'b11 &&
	     CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q4 ;
  assign NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1011_ETC___d371 =
	     { decoder_func_32_inst[6:2] != 5'b01011 &&
	       ((decoder_func_32_inst[6:2] == 5'b11000) ?
		  decoder_func_32_inst[7] :
		  decoder_func_32_inst[6:2] != 5'b01101 &&
		  decoder_func_32_inst[6:2] != 5'b00101 &&
		  ((decoder_func_32_inst[6:2] == 5'b11011) ?
		     decoder_func_32_inst[20] :
		     decoder_func_32_inst[31])),
	       CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q8,
	       CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q9,
	       decoder_func_32_inst[6:2] != 5'b01011 &&
	       ((decoder_func_32_inst[6:2] == 5'b01000) ?
		  decoder_func_32_inst[7] :
		  decoder_func_32_inst[6:2] != 5'b11000 &&
		  decoder_func_32_inst[6:2] != 5'b01101 &&
		  decoder_func_32_inst[6:2] != 5'b00101 &&
		  decoder_func_32_inst[6:2] != 5'b11011 &&
		  decoder_func_32_inst[20]) } ;
  assign _theResult_____6_snd__h1582 =
	     (decoder_func_32_inst[14:12] == 3'd0) ?
	       _theResult_____6_snd__h1609 :
	       6'd2 ;
  assign bit12_19__h46 = {8{decoder_func_32_inst[31]}} ;
  assign bit20_30__h47 =
	     { bit12_19__h46,
	       decoder_func_32_inst[31],
	       decoder_func_32_inst[31],
	       decoder_func_32_inst[31] } ;
  assign bit31__h48 =
	     decoder_func_32_inst[6:2] != 5'b01011 &&
	     decoder_func_32_inst[31] ;
  assign decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114 =
	     decoder_func_32_csrs[64] &&
	     (decoder_func_32_inst[14:12] == 3'd2 ||
	      decoder_func_32_inst[14:12] == 3'd3) &&
	     (decoder_func_32_inst[31:27] == 5'd0 ||
	      decoder_func_32_inst[31:27] == 5'd1 ||
	      decoder_func_32_inst[31:27] == 5'd3 ||
	      decoder_func_32_inst[31:27] == 5'd4 ||
	      decoder_func_32_inst[31:27] == 5'd8 ||
	      decoder_func_32_inst[31:27] == 5'd12 ||
	      decoder_func_32_inst[31:27] == 5'd16 ||
	      decoder_func_32_inst[31:27] == 5'd20 ||
	      decoder_func_32_inst[31:27] == 5'd24 ||
	      decoder_func_32_inst[31:27] == 5'd28 ||
	      decoder_func_32_inst[31:27] == 5'd2 &&
	      decoder_func_32_inst[24:20] == 5'd0) ;
  assign decoder_func_32_csrs_BIT_76_15_AND_decoder_fun_ETC___d127 =
	     decoder_func_32_csrs[76] &&
	     decoder_func_32_inst[31:25] == 7'd1 &&
	     (decoder_func_32_inst[14:12] == 3'd0 ||
	      !decoder_func_32_inst_BITS_14_TO_12_3_ULE_3___d121) ||
	     IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d126 ;
  assign decoder_func_32_inst_BITS_14_TO_12_3_ULE_3___d121 =
	     decoder_func_32_inst[14:12] <= 3'd3 ;
  assign decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84 =
	     decoder_func_32_inst[14:12] < 3'd4 ;
  assign decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158 =
	     decoder_func_32_inst[31:20] == 12'h002 &&
	     decoder_func_32_inst[19:15] == 5'd0 &&
	     decoder_func_32_inst[11:7] == 5'd0 &&
	     decoder_func_32_csrs[77] ||
	     decoder_func_32_inst[31:20] == 12'h302 &&
	     decoder_func_32_inst[19:15] == 5'd0 &&
	     decoder_func_32_inst[11:7] == 5'd0 &&
	     decoder_func_32_csrs[151:150] == 2'd3 ;
  assign decoder_func_32_inst_BIT_27_21_OR_decoder_func_ETC___d423 =
	     decoder_func_32_inst[27] | decoder_func_32_inst[28] ;
  assign fn___1__h4927 = { 3'd1, decoder_func_32_inst[12] } ;
  assign fn___1__h4949 = { 1'b1, decoder_func_32_inst[14:12] } ;
  assign immediate_value___1__h2154 =
	     { 15'd0,
	       decoder_func_32_inst[19:15],
	       NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1011_ETC___d371 } ;
  assign immediate_value__h49 =
	     { bit31__h48,
	       CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q10,
	       CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q11,
	       NOT_decoder_func_32_inst_BITS_6_TO_2_EQ_0b1011_ETC___d371 } ;
  assign instr_meta_funct__h352 =
	     (NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0b11_ETC___d192 ||
	      IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337) ?
	       temp1___1__h4863 :
	       temp1__h70 ;
  assign instr_meta_immediate__h351 =
	     ((decoder_func_32_inst[1:0] == 2'b11 ||
	       IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337) &&
	      decoder_func_32_inst[6:5] == 2'b11 &&
	      decoder_func_32_inst[4:2] == 3'b100 &&
	      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d340) ?
	       immediate_value___1__h2154 :
	       immediate_value__h49 ;
  assign temp1___1__h4863 = { 1'd0, x__h4866 } ;
  assign temp1__h70 =
	     { IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432,
	       decoder_func_32_inst[14:12] } ;
  assign trapcause___1__h1604 =
	     (decoder_func_32_csrs[84] &&
	      decoder_func_32_csrs[151:150] != 2'd3) ?
	       6'd8 :
	       6'd11 ;
  assign x__h194 =
	     (decoder_func_32_inst[6:2] == 5'b00100 ||
	      decoder_func_32_inst[6:2] == 5'b00110 ||
	      decoder_func_32_inst[6:2] == 5'b11100 ||
	      decoder_func_32_inst[6:2] == 5'b01101 ||
	      decoder_func_32_inst[6:2] == 5'b00101 ||
	      decoder_func_32_inst[6:2] == 5'b11011 ||
	      decoder_func_32_inst[6:2] == 5'b11001 ||
	      decoder_func_32_inst[6:4] == 3'b0) ?
	       5'd0 :
	       decoder_func_32_inst[24:20] ;
  assign x__h21 =
	     (decoder_func_32_inst[6:2] == 5'b01101 ||
	      decoder_func_32_inst[6:2] == 5'b00101 ||
	      decoder_func_32_inst[6:2] == 5'b11011 ||
	      decoder_func_32_inst[6:2] == 5'b11100 &&
	      decoder_func_32_inst[14]) ?
	       5'd0 :
	       decoder_func_32_inst[19:15] ;
  assign x__h4866 =
	     (NOT_decoder_func_32_inst_BITS_1_TO_0_6_EQ_0b11_ETC___d192 ||
	      decoder_func_32_inst[6:5] == 2'b0 ||
	      decoder_func_32_inst[6:5] == 2'b01) ?
	       6'd2 :
	       ((decoder_func_32_inst[6:5] == 2'b11) ?
		  _theResult_____6_snd__h1554 :
		  6'd2) ;
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[6:2])
      5'b01000, 5'b11000: x__h268 = 5'd0;
      default: x__h268 = decoder_func_32_inst[11:7];
    endcase
  end
  always@(decoder_func_32_inst or trapcause___1__h1604)
  begin
    case (decoder_func_32_inst[31:7])
      25'd0: _theResult_____6_snd__h1609 = trapcause___1__h1604;
      25'h0002000: _theResult_____6_snd__h1609 = 6'd3;
      default: _theResult_____6_snd__h1609 = 6'd2;
    endcase
  end
  always@(decoder_func_32_inst or _theResult_____6_snd__h1582)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0, 3'b001, 3'b011: _theResult_____6_snd__h1554 = 6'd2;
      3'b100: _theResult_____6_snd__h1554 = _theResult_____6_snd__h1582;
      default: _theResult_____6_snd__h1554 = 6'd2;
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[14:12])
      3'd0, 3'd5:
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119 =
	      decoder_func_32_inst[31:25] == 7'b0 ||
	      decoder_func_32_inst[31:25] == 7'b0100000;
      default: IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119 =
		   decoder_func_32_inst[31:25] == 7'b0;
    endcase
  end
  always@(decoder_func_32_inst or
	  decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158 or
	  decoder_func_32_csrs)
  begin
    case (decoder_func_32_inst[31:7])
      25'd0, 25'h0002000:
	  CASE_decoder_func_32_inst_BITS_31_TO_7_0_6_0x2_ETC__q1 = 4'd6;
      default: CASE_decoder_func_32_inst_BITS_31_TO_7_0_6_0x2_ETC__q1 =
		   decoder_func_32_inst_BITS_31_TO_20_44_EQ_0x2_4_ETC___d158 ?
		     4'd5 :
		     ((decoder_func_32_inst[31:20] == 12'h105 &&
		       decoder_func_32_inst[19:15] == 5'd0 &&
		       decoder_func_32_inst[11:7] == 5'd0 &&
		       decoder_func_32_csrs[151:150] == 2'd3) ?
			4'd7 :
			4'd6);
    endcase
  end
  always@(decoder_func_32_inst or
	  decoder_func_32_csrs_BIT_76_15_AND_decoder_fun_ETC___d127 or
	  decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84 or
	  decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114 or
	  decoder_func_32_csrs or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132 =
	      decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84;
      3'b011:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132 =
	      decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114;
      3'b100:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132 =
	      decoder_func_32_csrs[76] &&
	      decoder_func_32_inst[31:25] == 7'd1 ||
	      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d119;
      default: IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132 =
		   decoder_func_32_inst[4:2] == 3'b101 ||
		   decoder_func_32_inst[4:2] == 3'b110 &&
		   decoder_func_32_csrs_BIT_76_15_AND_decoder_fun_ETC___d127;
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d184)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2 =
	      decoder_func_32_inst[14:12] != 3'd2 &&
	      decoder_func_32_inst[14:12] != 3'd3;
      3'b001:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2 =
	      decoder_func_32_inst[14:12] == 3'd0;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2 =
		   decoder_func_32_inst[4:2] == 3'b011 ||
		   decoder_func_32_inst[4:2] == 3'b100 &&
		   IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d184;
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3 =
	      decoder_func_32_inst[14:12] != 3'd7;
      3'b011:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3 =
	      decoder_func_32_inst[14:12] == 3'd0 ||
	      decoder_func_32_inst[14:12] == 3'd1;
      3'b100:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3 =
	      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3 =
		   decoder_func_32_inst[4:2] == 3'b101 ||
		   decoder_func_32_inst[4:2] == 3'b110 &&
		   (decoder_func_32_inst[14:12] == 3'd0 ||
		    ((decoder_func_32_inst[14:12] == 3'd1) ?
		       decoder_func_32_inst[31:25] == 7'b0 :
		       decoder_func_32_inst[14:12] == 3'd5 &&
		       (decoder_func_32_inst[31:25] == 7'b0 ||
			decoder_func_32_inst[31:25] == 7'b0100000)));
    endcase
  end
  always@(decoder_func_32_inst or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2 or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3 or
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132)
  begin
    case (decoder_func_32_inst[6:5])
      2'b0:
	  CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q4 =
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q3;
      2'b01:
	  CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q4 =
	      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d132;
      default: CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q4 =
		   decoder_func_32_inst[6:5] == 2'b11 &&
		   CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_NOT__ETC__q2;
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[14:12])
      3'd0, 3'd5:
	  CASE_decoder_func_32_inst_BITS_14_TO_12_0_NOT__ETC__q5 =
	      decoder_func_32_inst[31:25] != 7'b0 &&
	      decoder_func_32_inst[31:25] != 7'b0100000;
      default: CASE_decoder_func_32_inst_BITS_14_TO_12_0_NOT__ETC__q5 =
		   decoder_func_32_inst[31:25] != 7'b0;
    endcase
  end
  always@(decoder_func_32_inst or
	  NOT_decoder_func_32_csrs_BIT_76_15_86_OR_NOT_d_ETC___d296 or
	  decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84 or
	  decoder_func_32_csrs or
	  CASE_decoder_func_32_inst_BITS_14_TO_12_0_NOT__ETC__q5)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301 =
	      !decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84;
      3'b011:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301 =
	      !decoder_func_32_csrs[64] ||
	      decoder_func_32_inst[14:12] != 3'd2 &&
	      decoder_func_32_inst[14:12] != 3'd3 ||
	      decoder_func_32_inst[31:27] != 5'd0 &&
	      decoder_func_32_inst[31:27] != 5'd1 &&
	      decoder_func_32_inst[31:27] != 5'd3 &&
	      decoder_func_32_inst[31:27] != 5'd4 &&
	      decoder_func_32_inst[31:27] != 5'd8 &&
	      decoder_func_32_inst[31:27] != 5'd12 &&
	      decoder_func_32_inst[31:27] != 5'd16 &&
	      decoder_func_32_inst[31:27] != 5'd20 &&
	      decoder_func_32_inst[31:27] != 5'd24 &&
	      decoder_func_32_inst[31:27] != 5'd28 &&
	      (decoder_func_32_inst[31:27] != 5'd2 ||
	       decoder_func_32_inst[24:20] != 5'd0);
      3'b100:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301 =
	      (!decoder_func_32_csrs[76] ||
	       decoder_func_32_inst[31:25] != 7'd1) &&
	      CASE_decoder_func_32_inst_BITS_14_TO_12_0_NOT__ETC__q5;
      default: IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301 =
		   decoder_func_32_inst[4:2] != 3'b101 &&
		   (decoder_func_32_inst[4:2] != 3'b110 ||
		    NOT_decoder_func_32_csrs_BIT_76_15_86_OR_NOT_d_ETC___d296);
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d330)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6 =
	      decoder_func_32_inst[14:12] == 3'd2 ||
	      decoder_func_32_inst[14:12] == 3'd3;
      3'b001:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6 =
	      decoder_func_32_inst[14:12] != 3'd0;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6 =
		   decoder_func_32_inst[4:2] != 3'b011 &&
		   (decoder_func_32_inst[4:2] != 3'b100 ||
		    IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d330);
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7 =
	      decoder_func_32_inst[14:12] == 3'd7;
      3'b011:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7 =
	      decoder_func_32_inst[14:12] != 3'd0 &&
	      decoder_func_32_inst[14:12] != 3'd1;
      3'b100:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7 =
	      (decoder_func_32_inst[14:12] == 3'd1) ?
		decoder_func_32_inst[31:26] != 6'd0 :
		decoder_func_32_inst[14:12] == 3'd5 &&
		decoder_func_32_inst[31:26] != 6'd0 &&
		decoder_func_32_inst[31:26] != 6'b010000;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7 =
		   decoder_func_32_inst[4:2] != 3'b101 &&
		   (decoder_func_32_inst[4:2] != 3'b110 ||
		    decoder_func_32_inst[14:12] != 3'd0 &&
		    ((decoder_func_32_inst[14:12] == 3'd1) ?
		       decoder_func_32_inst[31:25] != 7'b0 :
		       decoder_func_32_inst[14:12] != 3'd5 ||
		       decoder_func_32_inst[31:25] != 7'b0 &&
		       decoder_func_32_inst[31:25] != 7'b0100000));
    endcase
  end
  always@(decoder_func_32_inst or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6 or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7 or
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301)
  begin
    case (decoder_func_32_inst[6:5])
      2'b0:
	  IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337 =
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q7;
      2'b01:
	  IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337 =
	      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d301;
      default: IF_decoder_func_32_inst_BITS_6_TO_5_9_EQ_0b0_0_ETC___d337 =
		   decoder_func_32_inst[6:5] != 2'b11 ||
		   CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_deco_ETC__q6;
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00101, 5'b01011, 5'b01101:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q8 = 6'd0;
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q8 =
		   decoder_func_32_inst[30:25];
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00101, 5'b01011, 5'b01101:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q9 = 4'd0;
      5'b01000, 5'b11000:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q9 =
	      decoder_func_32_inst[11:8];
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_0__ETC__q9 =
		   decoder_func_32_inst[24:21];
    endcase
  end
  always@(decoder_func_32_inst or bit20_30__h47)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00101, 5'b01101:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q10 =
	      decoder_func_32_inst[30:20];
      5'b01011:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q10 = 11'd0;
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q10 =
		   bit20_30__h47;
    endcase
  end
  always@(decoder_func_32_inst or bit12_19__h46)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00101, 5'b01101, 5'b11011:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q11 =
	      decoder_func_32_inst[19:12];
      5'b01011:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q11 = 8'd0;
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b101_de_ETC__q11 =
		   bit12_19__h46;
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411)
  begin
    case (decoder_func_32_inst[14:12])
      3'd2: fn___1__h4966 = 4'b1100;
      3'd3: fn___1__h4966 = 4'b1110;
      3'd5:
	  fn___1__h4966 =
	      IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411;
      default: fn___1__h4966 = { 1'b0, decoder_func_32_inst[14:12] };
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411)
  begin
    case (decoder_func_32_inst[14:12])
      3'd0: fn___1__h5028 = decoder_func_32_inst[30] ? 4'b1010 : 4'b0;
      3'd2: fn___1__h5028 = 4'b1100;
      3'd3: fn___1__h5028 = 4'b1110;
      3'd5:
	  fn___1__h5028 =
	      IF_decoder_func_32_inst_BIT_30_10_THEN_0b1011__ETC___d411;
      default: fn___1__h5028 = { 1'b0, decoder_func_32_inst[14:12] };
    endcase
  end
  always@(decoder_func_32_inst or
	  fn___1__h4966 or
	  decoder_func_32_inst_BIT_27_21_OR_decoder_func_ETC___d423 or
	  fn___1__h5028 or fn___1__h4949 or fn___1__h4927)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00100, 5'b00110:
	  IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432 =
	      fn___1__h4966;
      5'b01011:
	  IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432 =
	      { decoder_func_32_inst_BIT_27_21_OR_decoder_func_ETC___d423 ?
		  decoder_func_32_inst[29:27] :
		  decoder_func_32_inst[31:29],
		decoder_func_32_inst_BIT_27_21_OR_decoder_func_ETC___d423 ||
		decoder_func_32_inst[27] };
      5'b01100, 5'b01110:
	  IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432 =
	      fn___1__h5028;
      5'b11000:
	  IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432 =
	      decoder_func_32_inst[14] ? fn___1__h4949 : fn___1__h4927;
      default: IF_decoder_func_32_inst_BITS_6_TO_2_EQ_0b11000_ETC___d432 =
		   4'd0;
    endcase
  end
  always@(decoder_func_32_inst or
	  decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84 or
	  decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114 or
	  IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d205 or
	  IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d207)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 =
	      decoder_func_32_inst_BITS_14_TO_12_3_ULT_4___d84 ? 4'd1 : 4'd6;
      3'b011:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 =
	      decoder_func_32_csrs_BIT_64_5_AND_decoder_func_ETC___d114 ?
		4'd1 :
		4'd6;
      3'b100:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 =
	      IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d205;
      3'b101:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 = 4'd0;
      3'b110:
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 =
	      IF_decoder_func_32_csrs_BIT_76_15_AND_decoder__ETC___d207;
      default: IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 =
		   4'd6;
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[14:12])
      3'd0, 3'd1:
	  CASE_decoder_func_32_inst_BITS_14_TO_12_0_1_1_1_6__q12 = 4'd1;
      default: CASE_decoder_func_32_inst_BITS_14_TO_12_0_1_1_1_6__q12 = 4'd6;
    endcase
  end
  always@(decoder_func_32_inst or
	  CASE_decoder_func_32_inst_BITS_14_TO_12_0_1_1_1_6__q12 or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 =
	      (decoder_func_32_inst[14:12] == 3'd7) ? 4'd6 : 4'd1;
      3'b011:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 =
	      CASE_decoder_func_32_inst_BITS_14_TO_12_0_1_1_1_6__q12;
      3'b100:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 =
	      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_1_8_ETC___d68 ?
		4'd0 :
		4'd6;
      3'b101: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 = 4'd0;
      3'b110:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 =
	      (decoder_func_32_inst[14:12] == 3'd0 ||
	       ((decoder_func_32_inst[14:12] == 3'd1) ?
		  decoder_func_32_inst[31:25] == 7'b0 :
		  decoder_func_32_inst[14:12] == 3'd5 &&
		  (decoder_func_32_inst[31:25] == 7'b0 ||
		   decoder_func_32_inst[31:25] == 7'b0100000))) ?
		4'd0 :
		4'd6;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 = 4'd6;
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d220)
  begin
    case (decoder_func_32_inst[4:2])
      3'b0:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14 =
	      (decoder_func_32_inst[14:12] != 3'd2 &&
	       decoder_func_32_inst[14:12] != 3'd3) ?
		4'd2 :
		4'd6;
      3'b001:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14 =
	      (decoder_func_32_inst[14:12] == 3'd0) ? 4'd4 : 4'd6;
      3'b011: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14 = 4'd3;
      3'b100:
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14 =
	      IF_decoder_func_32_inst_BITS_14_TO_12_3_EQ_0_7_ETC___d220;
      default: CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14 = 4'd6;
    endcase
  end
  always@(decoder_func_32_inst or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13 or
	  IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212 or
	  CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14)
  begin
    case (decoder_func_32_inst[6:5])
      2'b0:
	  CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15 =
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_d_ETC__q13;
      2'b01:
	  CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15 =
	      IF_decoder_func_32_inst_BITS_4_TO_2_1_EQ_0b0_2_ETC___d212;
      2'd2: CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15 = 4'd6;
      2'b11:
	  CASE_decoder_func_32_inst_BITS_6_TO_5_0b0_CASE_ETC__q15 =
	      CASE_decoder_func_32_inst_BITS_4_TO_2_0b0_IF_N_ETC__q14;
    endcase
  end
  always@(decoder_func_32_inst)
  begin
    case (decoder_func_32_inst[6:2])
      5'b00011:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b11_3_0_ETC__q16 = 2'd3;
      5'b01000:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b11_3_0_ETC__q16 = 2'd1;
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b11_3_0_ETC__q16 = 2'd2;
    endcase
  end
  always@(decoder_func_32_inst or
	  IF_decoder_func_32_compressed_THEN_3_ELSE_2___d40)
  begin
    case (decoder_func_32_inst[6:2])
      5'b0, 5'b00100, 5'b00101, 5'b00110, 5'b01101:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b0_1_0b_ETC__q17 = 2'd1;
      5'b00011, 5'b11001, 5'b11011:
	  CASE_decoder_func_32_inst_BITS_6_TO_2_0b0_1_0b_ETC__q17 =
	      IF_decoder_func_32_compressed_THEN_3_ELSE_2___d40;
      default: CASE_decoder_func_32_inst_BITS_6_TO_2_0b0_1_0b_ETC__q17 = 2'd0;
    endcase
  end
endmodule  // module_decoder_func_32

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:53 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// decode_word32                  O     1
// decode_word32_inst             I    32
// decode_word32_misa_c           I     1
//
// Combinational paths from inputs to outputs:
//   (decode_word32_inst, decode_word32_misa_c) -> decode_word32
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_decode_word32(decode_word32_inst,
			    decode_word32_misa_c,
			    decode_word32);
  // value method decode_word32
  input  [31 : 0] decode_word32_inst;
  input  decode_word32_misa_c;
  output decode_word32;

  // signals for module outputs
  wire decode_word32;

  // value method decode_word32
  assign decode_word32 =
	     (decode_word32_misa_c && decode_word32_inst[1:0] != 2'b11) ?
	       decode_word32_inst[1:0] == 2'd1 &&
	       (decode_word32_inst[15:13] == 3'b001 ||
		decode_word32_inst[15:13] == 3'b100 &&
		decode_word32_inst[12:10] == 3'b111 &&
		!decode_word32_inst[6]) :
	       decode_word32_inst[6:2] == 5'b00110 ||
	       decode_word32_inst[6:2] == 5'b01110 ||
	       decode_word32_inst[6:3] == 4'b0101 && !decode_word32_inst[12] ;
endmodule  // module_decode_word32

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:13 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// fn_alu                         O   138
// fn_alu_fn                      I     4
// fn_alu_op1                     I    64
// fn_alu_op2                     I    64
// fn_alu_op3                     I    64
// fn_alu_imm_value               I    64
// fn_alu_inst_type               I     4
// fn_alu_funct3                  I     3
// fn_alu_memaccess               I     2
// fn_alu_word32                  I     1
// fn_alu_misa_c                  I     1
// fn_alu_lpc                     I     2 unused
// fn_alu_tdata1                  I    44
// fn_alu_tdata2                  I   128
// fn_alu_tenable                 I     2
//
// Combinational paths from inputs to outputs:
//   (fn_alu_fn,
//    fn_alu_op1,
//    fn_alu_op2,
//    fn_alu_op3,
//    fn_alu_imm_value,
//    fn_alu_inst_type,
//    fn_alu_funct3,
//    fn_alu_memaccess,
//    fn_alu_word32,
//    fn_alu_misa_c,
//    fn_alu_tdata1,
//    fn_alu_tdata2,
//    fn_alu_tenable) -> fn_alu
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_fn_alu(fn_alu_fn,
		     fn_alu_op1,
		     fn_alu_op2,
		     fn_alu_op3,
		     fn_alu_imm_value,
		     fn_alu_inst_type,
		     fn_alu_funct3,
		     fn_alu_memaccess,
		     fn_alu_word32,
		     fn_alu_misa_c,
		     fn_alu_lpc,
		     fn_alu_tdata1,
		     fn_alu_tdata2,
		     fn_alu_tenable,
		     fn_alu);
  // value method fn_alu
  input  [3 : 0] fn_alu_fn;
  input  [63 : 0] fn_alu_op1;
  input  [63 : 0] fn_alu_op2;
  input  [63 : 0] fn_alu_op3;
  input  [63 : 0] fn_alu_imm_value;
  input  [3 : 0] fn_alu_inst_type;
  input  [2 : 0] fn_alu_funct3;
  input  [1 : 0] fn_alu_memaccess;
  input  fn_alu_word32;
  input  fn_alu_misa_c;
  input  [1 : 0] fn_alu_lpc;
  input  [43 : 0] fn_alu_tdata1;
  input  [127 : 0] fn_alu_tdata2;
  input  [1 : 0] fn_alu_tenable;
  output [137 : 0] fn_alu;

  // signals for module outputs
  wire [137 : 0] fn_alu;

  // remaining internal signals
  reg [63 : 0] final_output__h57, shin__h53;
  reg [1 : 0] CASE_fn_alu_inst_type_1_0_5_1_2__q5;
  reg CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2,
      CASE_fn_alu_tdata1_BITS_14_TO_11_2_IF_fn_alu_t_ETC__q1,
      IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97,
      IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144,
      IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147;
  wire [64 : 0] fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371,
		fn_alu_fn_BIT_3_AND_shin3_BIT_63_CONCAT_shin3__q3,
		inv_op2__h41,
		x__h2126;
  wire [63 : 0] _theResult_____7__h59,
		_theResult____h1546,
		_theResult____h876,
		effective_address__h58,
		final_output___1__h2086,
		op1_xor_op2__h42,
		result__h942,
		shift_inright__h52,
		shift_l__h56,
		x__h2082;
  wire [31 : 0] final_output7_BITS_31_TO_0__q4, upper_bits__h51;
  wire [6 : 0] IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d495;
  wire [5 : 0] _theResult_____4_fst__h1839,
	       _theResult_____5_fst__h1870,
	       cause___1__h1841,
	       cause___1__h1886,
	       cause__h60,
	       cause__h63,
	       cause__h66,
	       shift_amt__h50;
  wire [1 : 0] IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d209;
  wire IF_NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu__ETC___d203,
       IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61,
       IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d96,
       IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132,
       INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190,
       NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu_ins_ETC___d165,
       NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49,
       NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142,
       NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d71,
       adder_z_flag__h44,
       fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_BI_ETC___d149,
       fn_alu_inst_type_EQ_2_72_AND_IF_fn_alu_fn_EQ_2_ETC___d195,
       fn_alu_inst_type_EQ_4_4_OR_fn_alu_inst_type_EQ_ETC___d200,
       fn_alu_tdata1_BIT_19_AND_fn_alu_memaccess_EQ_0_ETC___d89,
       fn_alu_tdata1_BIT_41_02_AND_fn_alu_memaccess_E_ETC___d124,
       fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140,
       fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66,
       fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138,
       fn_alu_tenable_BIT_1_AND_NOT_fn_alu_tenable_BI_ETC___d127,
       sign__h45,
       x__h10053;

  // value method fn_alu
  assign fn_alu =
	     { 1'd1,
	       IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d209,
	       x__h2082,
	       _theResult_____7__h59,
	       IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d495 } ;

  // remaining internal signals
  assign IF_NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu__ETC___d203 =
	     (fn_alu_memaccess != 2'd3 && fn_alu_inst_type == 4'd1) ?
	       _theResult_____7__h59[63:32] != 32'd0 :
	       fn_alu_inst_type_EQ_4_4_OR_fn_alu_inst_type_EQ_ETC___d200 ||
	       fn_alu_inst_type == 4'd6 ;
  assign IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d209 =
	     (fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_BI_ETC___d149 ||
	      NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu_ins_ETC___d165 ||
	      IF_NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu__ETC___d203) ?
	       2'd3 :
	       CASE_fn_alu_inst_type_1_0_5_1_2__q5 ;
  assign IF_fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_ETC___d495 =
	     { fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_BI_ETC___d149 ?
		 6'd3 :
		 _theResult_____4_fst__h1839,
	       fn_alu_inst_type_EQ_2_72_AND_IF_fn_alu_fn_EQ_2_ETC___d195 ||
	       fn_alu_inst_type == 4'd4 ||
	       fn_alu_inst_type == 4'd3 } ;
  assign IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61 =
	     _theResult____h876 < fn_alu_tdata2[63:0] ;
  assign IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d96 =
	     IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61 ||
	     ((fn_alu_tdata1[14:11] == 4'd2) ?
		!IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61 :
		fn_alu_tdata1[14:11] == 4'd0 &&
		fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66) ;
  assign IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 =
	     _theResult____h1546 < fn_alu_tdata2[127:64] ;
  assign INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190 =
	     ({ sign__h45 & fn_alu_op1[63], fn_alu_op1 } ^
	      65'h10000000000000000) <
	     ({ sign__h45 & fn_alu_op2[63], fn_alu_op2 } ^
	      65'h10000000000000000) ;
  assign NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu_ins_ETC___d165 =
	     fn_alu_memaccess != 2'd3 && fn_alu_inst_type == 4'd1 &&
	     (fn_alu_funct3[1:0] == 2'd1 && effective_address__h58[0] ||
	      fn_alu_funct3[1:0] == 2'd2 &&
	      _theResult_____7__h59[1:0] != 2'd0 ||
	      fn_alu_funct3[1:0] == 2'd3 &&
	      effective_address__h58[2:0] != 3'd0) ;
  assign NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 =
	     (!fn_alu_tdata1[19] || fn_alu_memaccess != 2'd0 ||
	      fn_alu_tdata1[1]) &&
	     (!fn_alu_tdata1[18] || fn_alu_memaccess != 2'd1) ||
	     fn_alu_tdata1[5:2] != 4'd0 &&
	     (fn_alu_tdata1[5:2] != 4'd1 || fn_alu_funct3[1:0] != 2'd0) &&
	     (fn_alu_tdata1[5:2] != 4'd2 || fn_alu_funct3[1:0] != 2'd1) &&
	     (fn_alu_tdata1[5:2] != 4'd3 || fn_alu_funct3[1:0] != 2'd2) &&
	     (fn_alu_tdata1[5:2] != 4'd5 || fn_alu_funct3[1:0] != 2'd3) ;
  assign NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142 =
	     (!fn_alu_tenable[0] || fn_alu_tdata1[21:20] != 2'd0 ||
	      NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 ||
	      !fn_alu_tdata1[10]) &&
	     ((fn_alu_tdata1[36:33] == 4'd0) ?
		fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140 :
		fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138) ;
  assign NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d71 =
	     !fn_alu_tenable[0] || fn_alu_tdata1[21:20] != 2'd0 ||
	     NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 ||
	     CASE_fn_alu_tdata1_BITS_14_TO_11_2_IF_fn_alu_t_ETC__q1 ;
  assign _theResult_____4_fst__h1839 =
	     NOT_fn_alu_memaccess_EQ_3_50_51_AND_fn_alu_ins_ETC___d165 ?
	       cause___1__h1841 :
	       cause__h66 ;
  assign _theResult_____5_fst__h1870 =
	     (_theResult_____7__h59[63:32] == 32'd0) ?
	       cause__h63 :
	       cause___1__h1886 ;
  assign _theResult_____7__h59 =
	     (fn_alu_inst_type == 4'd4) ?
	       result__h942 :
	       effective_address__h58 ;
  assign _theResult____h1546 =
	     fn_alu_tdata1[23] ? fn_alu_op2 : _theResult_____7__h59 ;
  assign _theResult____h876 =
	     fn_alu_tdata1[1] ? fn_alu_op2 : _theResult_____7__h59 ;
  assign adder_z_flag__h44 = ~(op1_xor_op2__h42 != 64'd0) ;
  assign cause___1__h1841 = (fn_alu_memaccess == 2'd0) ? cause__h66 : 6'd6 ;
  assign cause___1__h1886 = (fn_alu_memaccess == 2'd0) ? 6'd5 : 6'd7 ;
  assign cause__h60 =
	     (fn_alu_inst_type == 4'd6) ?
	       { fn_alu_fn[2:0], fn_alu_funct3 } :
	       6'd4 ;
  assign cause__h63 =
	     fn_alu_inst_type_EQ_4_4_OR_fn_alu_inst_type_EQ_ETC___d200 ?
	       6'd0 :
	       cause__h60 ;
  assign cause__h66 =
	     (fn_alu_memaccess != 2'd3 && fn_alu_inst_type == 4'd1) ?
	       _theResult_____5_fst__h1870 :
	       cause__h63 ;
  assign effective_address__h58 = fn_alu_op3 + fn_alu_imm_value ;
  assign final_output7_BITS_31_TO_0__q4 = final_output__h57[31:0] ;
  assign final_output___1__h2086 =
	     { {32{final_output7_BITS_31_TO_0__q4[31]}},
	       final_output7_BITS_31_TO_0__q4 } ;
  assign fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371 =
	     { fn_alu_fn[3] & shin__h53[63], shin__h53 } >> shift_amt__h50 |
	     ~(65'h1FFFFFFFFFFFFFFFF >> shift_amt__h50) &
	     {65{fn_alu_fn_BIT_3_AND_shin3_BIT_63_CONCAT_shin3__q3[64]}} ;
  assign fn_alu_fn_BIT_3_AND_shin3_BIT_63_CONCAT_shin3__q3 =
	     { fn_alu_fn[3] & shin__h53[63], shin__h53 } ;
  assign fn_alu_inst_type_EQ_1_AND_IF_fn_alu_tenable_BI_ETC___d149 =
	     fn_alu_inst_type == 4'd1 &&
	     (fn_alu_tenable_BIT_1_AND_NOT_fn_alu_tenable_BI_ETC___d127 ?
		IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147 :
		fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138) ;
  assign fn_alu_inst_type_EQ_2_72_AND_IF_fn_alu_fn_EQ_2_ETC___d195 =
	     fn_alu_inst_type == 4'd2 &&
	     CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2 ;
  assign fn_alu_inst_type_EQ_4_4_OR_fn_alu_inst_type_EQ_ETC___d200 =
	     (fn_alu_inst_type == 4'd4 || fn_alu_inst_type == 4'd3 ||
	      fn_alu_inst_type_EQ_2_72_AND_IF_fn_alu_fn_EQ_2_ETC___d195) &&
	     _theResult_____7__h59[1] &&
	     !fn_alu_misa_c ;
  assign fn_alu_tdata1_BIT_19_AND_fn_alu_memaccess_EQ_0_ETC___d89 =
	     (fn_alu_tdata1[19] && fn_alu_memaccess == 2'd0 &&
	      !fn_alu_tdata1[1] ||
	      fn_alu_tdata1[18] && fn_alu_memaccess == 2'd1) &&
	     (fn_alu_tdata1[5:2] == 4'd0 ||
	      fn_alu_tdata1[5:2] == 4'd1 && fn_alu_funct3[1:0] == 2'd0 ||
	      fn_alu_tdata1[5:2] == 4'd2 && fn_alu_funct3[1:0] == 2'd1 ||
	      fn_alu_tdata1[5:2] == 4'd3 && fn_alu_funct3[1:0] == 2'd2 ||
	      fn_alu_tdata1[5:2] == 4'd5 && fn_alu_funct3[1:0] == 2'd3) ;
  assign fn_alu_tdata1_BIT_41_02_AND_fn_alu_memaccess_E_ETC___d124 =
	     (fn_alu_tdata1[41] && fn_alu_memaccess == 2'd0 &&
	      !fn_alu_tdata1[23] ||
	      fn_alu_tdata1[40] && fn_alu_memaccess == 2'd1) &&
	     (fn_alu_tdata1[27:24] == 4'd0 ||
	      fn_alu_tdata1[27:24] == 4'd1 && fn_alu_funct3[1:0] == 2'd0 ||
	      fn_alu_tdata1[27:24] == 4'd2 && fn_alu_funct3[1:0] == 2'd1 ||
	      fn_alu_tdata1[27:24] == 4'd3 && fn_alu_funct3[1:0] == 2'd2 ||
	      fn_alu_tdata1[27:24] == 4'd5 && fn_alu_funct3[1:0] == 2'd3) ;
  assign fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140 =
	     fn_alu_tdata2[127:64] == _theResult____h1546 ||
	     !fn_alu_tdata1[10] &&
	     fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138 ;
  assign fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66 =
	     fn_alu_tdata2[63:0] == _theResult____h876 ;
  assign fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138 =
	     fn_alu_tenable[0] && fn_alu_tdata1[21:20] == 2'd0 &&
	     fn_alu_tdata1_BIT_19_AND_fn_alu_memaccess_EQ_0_ETC___d89 &&
	     IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97 ;
  assign fn_alu_tenable_BIT_1_AND_NOT_fn_alu_tenable_BI_ETC___d127 =
	     fn_alu_tenable[1] &&
	     (NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d71 &&
	      (!fn_alu_tenable[0] || fn_alu_tdata1[21:20] != 2'd0 ||
	       NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 ||
	       !fn_alu_tdata1[10]) ||
	      fn_alu_tenable[0] && fn_alu_tdata1[21:20] == 2'd0 &&
	      fn_alu_tdata1_BIT_19_AND_fn_alu_memaccess_EQ_0_ETC___d89 &&
	      fn_alu_tdata1[10] &&
	      IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97) &&
	     fn_alu_tdata1[43:42] == 2'd0 &&
	     fn_alu_tdata1_BIT_41_02_AND_fn_alu_memaccess_E_ETC___d124 ;
  assign inv_op2__h41 = { fn_alu_op2 ^ {64{fn_alu_fn[1]}}, fn_alu_fn[1] } ;
  assign op1_xor_op2__h42 = fn_alu_op1 ^ fn_alu_op2 ;
  assign result__h942 = { effective_address__h58[63:1], 1'd0 } ;
  assign shift_amt__h50 =
	     { !fn_alu_word32 && fn_alu_op2[5], fn_alu_op2[4:0] } ;
  assign shift_inright__h52 = { upper_bits__h51, fn_alu_op1[31:0] } ;
  assign shift_l__h56 =
	     { fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[0],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[1],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[2],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[3],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[4],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[5],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[6],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[7],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[8],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[9],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[10],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[11],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[12],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[13],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[14],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[15],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[16],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[17],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[18],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[19],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[20],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[21],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[22],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[23],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[24],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[25],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[26],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[27],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[28],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[29],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[30],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[31],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[32],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[33],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[34],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[35],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[36],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[37],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[38],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[39],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[40],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[41],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[42],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[43],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[44],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[45],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[46],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[47],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[48],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[49],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[50],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[51],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[52],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[53],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[54],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[55],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[56],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[57],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[58],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[59],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[60],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[61],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[62],
	       fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[63] } ;
  assign sign__h45 = ~fn_alu_fn[1] ;
  assign upper_bits__h51 =
	     fn_alu_word32 ? {32{x__h10053}} : fn_alu_op1[63:32] ;
  assign x__h10053 = fn_alu_fn[3] & fn_alu_op1[31] ;
  assign x__h2082 =
	     fn_alu_word32 ? final_output___1__h2086 : final_output__h57 ;
  assign x__h2126 = { fn_alu_op1, 1'b1 } + inv_op2__h41 ;
  always@(fn_alu_fn or fn_alu_op1 or upper_bits__h51 or shift_inright__h52)
  begin
    case (fn_alu_fn)
      4'd5, 4'd11: shin__h53 = shift_inright__h52;
      default: shin__h53 =
		   { fn_alu_op1[0],
		     fn_alu_op1[1],
		     fn_alu_op1[2],
		     fn_alu_op1[3],
		     fn_alu_op1[4],
		     fn_alu_op1[5],
		     fn_alu_op1[6],
		     fn_alu_op1[7],
		     fn_alu_op1[8],
		     fn_alu_op1[9],
		     fn_alu_op1[10],
		     fn_alu_op1[11],
		     fn_alu_op1[12],
		     fn_alu_op1[13],
		     fn_alu_op1[14],
		     fn_alu_op1[15],
		     fn_alu_op1[16],
		     fn_alu_op1[17],
		     fn_alu_op1[18],
		     fn_alu_op1[19],
		     fn_alu_op1[20],
		     fn_alu_op1[21],
		     fn_alu_op1[22],
		     fn_alu_op1[23],
		     fn_alu_op1[24],
		     fn_alu_op1[25],
		     fn_alu_op1[26],
		     fn_alu_op1[27],
		     fn_alu_op1[28],
		     fn_alu_op1[29],
		     fn_alu_op1[30],
		     fn_alu_op1[31],
		     upper_bits__h51[0],
		     upper_bits__h51[1],
		     upper_bits__h51[2],
		     upper_bits__h51[3],
		     upper_bits__h51[4],
		     upper_bits__h51[5],
		     upper_bits__h51[6],
		     upper_bits__h51[7],
		     upper_bits__h51[8],
		     upper_bits__h51[9],
		     upper_bits__h51[10],
		     upper_bits__h51[11],
		     upper_bits__h51[12],
		     upper_bits__h51[13],
		     upper_bits__h51[14],
		     upper_bits__h51[15],
		     upper_bits__h51[16],
		     upper_bits__h51[17],
		     upper_bits__h51[18],
		     upper_bits__h51[19],
		     upper_bits__h51[20],
		     upper_bits__h51[21],
		     upper_bits__h51[22],
		     upper_bits__h51[23],
		     upper_bits__h51[24],
		     upper_bits__h51[25],
		     upper_bits__h51[26],
		     upper_bits__h51[27],
		     upper_bits__h51[28],
		     upper_bits__h51[29],
		     upper_bits__h51[30],
		     upper_bits__h51[31] };
    endcase
  end
  always@(fn_alu_tdata1 or
	  fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66 or
	  IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61)
  begin
    case (fn_alu_tdata1[14:11])
      4'd2:
	  CASE_fn_alu_tdata1_BITS_14_TO_11_2_IF_fn_alu_t_ETC__q1 =
	      IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61;
      4'd3:
	  CASE_fn_alu_tdata1_BITS_14_TO_11_2_IF_fn_alu_t_ETC__q1 =
	      !IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61;
      default: CASE_fn_alu_tdata1_BITS_14_TO_11_2_IF_fn_alu_t_ETC__q1 =
		   fn_alu_tdata1[14:11] != 4'd0 ||
		   !fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66;
    endcase
  end
  always@(fn_alu_tdata1 or
	  fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66 or
	  IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61 or
	  IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d96)
  begin
    case (fn_alu_tdata1[14:11])
      4'd2:
	  IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97 =
	      !IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d61;
      4'd3:
	  IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97 =
	      IF_fn_alu_tdata1_BIT_1_3_THEN_fn_alu_op2_ELSE__ETC___d96;
      default: IF_fn_alu_tdata1_BITS_14_TO_11_2_EQ_3_3_THEN_I_ETC___d97 =
		   fn_alu_tdata1[14:11] == 4'd0 &&
		   fn_alu_tdata2_BITS_63_TO_0_0_EQ_IF_fn_alu_tdat_ETC___d66;
    endcase
  end
  always@(fn_alu_tdata1 or
	  fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138 or
	  fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140 or
	  IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 or
	  NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142)
  begin
    case (fn_alu_tdata1[36:33])
      4'd0:
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144 =
	      fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140;
      4'd2:
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144 =
	      !IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 ||
	      NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142;
      default: IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144 =
		   fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138;
    endcase
  end
  always@(fn_alu_fn or
	  INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190 or
	  adder_z_flag__h44 or op1_xor_op2__h42)
  begin
    case (fn_alu_fn)
      4'd2:
	  CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2 =
	      adder_z_flag__h44;
      4'd3:
	  CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2 =
	      op1_xor_op2__h42 != 64'd0;
      4'd12, 4'd14:
	  CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2 =
	      INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190;
      default: CASE_fn_alu_fn_2_adder_z_flag4_3_NOT_op1_xor_o_ETC__q2 =
		   !INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190;
    endcase
  end
  always@(fn_alu_tdata1 or
	  fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138 or
	  fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140 or
	  IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 or
	  NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142 or
	  fn_alu_tenable or
	  NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 or
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144)
  begin
    case (fn_alu_tdata1[36:33])
      4'd0:
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147 =
	      fn_alu_tdata2_BITS_127_TO_64_31_EQ_IF_fn_alu_t_ETC___d140;
      4'd2:
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147 =
	      !IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 ||
	      NOT_fn_alu_tenable_BIT_0_OR_NOT_fn_alu_tdata1__ETC___d142;
      4'd3:
	  IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147 =
	      IF_fn_alu_tdata1_BIT_23_04_THEN_fn_alu_op2_ELS_ETC___d132 ||
	      (!fn_alu_tenable[0] || fn_alu_tdata1[21:20] != 2'd0 ||
	       NOT_fn_alu_tdata1_BIT_19_OR_NOT_fn_alu_memacce_ETC___d49 ||
	       !fn_alu_tdata1[10]) &&
	      IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_2_33_THEN_ETC___d144;
      default: IF_fn_alu_tdata1_BITS_36_TO_33_28_EQ_3_29_THEN_ETC___d147 =
		   fn_alu_tenable_BIT_0_AND_fn_alu_tdata1_BITS_21_ETC___d138;
    endcase
  end
  always@(fn_alu_fn or
	  op1_xor_op2__h42 or
	  x__h2126 or
	  shift_l__h56 or
	  fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371 or
	  fn_alu_op1 or
	  fn_alu_op2 or
	  INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190)
  begin
    case (fn_alu_fn)
      4'd0, 4'd10: final_output__h57 = x__h2126[64:1];
      4'd1: final_output__h57 = shift_l__h56;
      4'd5, 4'd11:
	  final_output__h57 =
	      fn_alu_fn_BIT_3_59_AND_IF_fn_alu_fn_EQ_5_56_OR_ETC___d371[63:0];
      4'd6: final_output__h57 = fn_alu_op1 | fn_alu_op2;
      4'd7: final_output__h57 = fn_alu_op1 & fn_alu_op2;
      4'd12, 4'd13, 4'd14, 4'd15:
	  final_output__h57 =
	      { 63'd0,
		INV_fn_alu_fn_BIT_1_82_83_AND_fn_alu_op1_BIT_6_ETC___d190 };
      default: final_output__h57 = op1_xor_op2__h42;
    endcase
  end
  always@(fn_alu_inst_type)
  begin
    case (fn_alu_inst_type)
      4'd1: CASE_fn_alu_inst_type_1_0_5_1_2__q5 = 2'd0;
      4'd5: CASE_fn_alu_inst_type_1_0_5_1_2__q5 = 2'd1;
      default: CASE_fn_alu_inst_type_1_0_5_1_2__q5 = 2'd2;
    endcase
  end
endmodule  // module_fn_alu

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:05 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// fn_decompress                  O    32
// fn_decompress_inst             I    16
//
// Combinational paths from inputs to outputs:
//   fn_decompress_inst -> fn_decompress
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_fn_decompress(fn_decompress_inst,
			    fn_decompress);
  // value method fn_decompress
  input  [15 : 0] fn_decompress_inst;
  output [31 : 0] fn_decompress;

  // signals for module outputs
  wire [31 : 0] fn_decompress;

  // remaining internal signals
  wire [31 : 0] IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d319,
		IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d322,
		IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1000__ETC___d321,
		IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1001__ETC___d318,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b100_8_ETC___d335,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b10_2__ETC___d324,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b110_8_ETC___d317,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b111_7_ETC___d343,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b11_2__ETC___d345,
		IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b1_2_A_ETC___d341,
		IF_fn_decompress_inst_BITS_15_TO_7_3_EQ_0b1110_ETC___d339;
  wire [11 : 0] SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67;
  wire [9 : 0] x__h1408, x__h4254;
  wire [8 : 0] x__h12235;
  wire [7 : 0] x__h12096, x__h1733;
  wire [6 : 0] x__h1569;
  wire [5 : 0] fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1;
  wire [3 : 0] x__h14618;
  wire [2 : 0] x__h14479, x__h2058;
  wire [1 : 0] x__h1873;
  wire fn_decompress_inst_BIT_10_AND_fn_decompress_in_ETC___d277,
       fn_decompress_inst_BIT_5_4_AND_fn_decompress_i_ETC___d288;

  // value method fn_decompress
  assign fn_decompress =
	     (fn_decompress_inst[15:12] == 4'b0001 &&
	      fn_decompress_inst[1:0] == 2'b0 ||
	      fn_decompress_inst[15:13] == 3'b0 &&
	      (fn_decompress_inst[11] || fn_decompress_inst[10] ||
	       fn_decompress_inst[9] ||
	       fn_decompress_inst[8] ||
	       fn_decompress_inst[7] ||
	       fn_decompress_inst[6] ||
	       fn_decompress_inst[5]) &&
	      fn_decompress_inst[1:0] == 2'b0) ?
	       { 2'd0, x__h1408, 10'd65, fn_decompress_inst[4:2], 7'd19 } :
	       ((fn_decompress_inst[15:13] == 3'b010 &&
		 fn_decompress_inst[1:0] == 2'b0) ?
		  { 5'd0,
		    x__h1569,
		    2'b01,
		    fn_decompress_inst[9:7],
		    5'b01001,
		    fn_decompress_inst[4:2],
		    7'd3 } :
		  IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b11_2__ETC___d345) ;

  // remaining internal signals
  assign IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d319 =
	     (fn_decompress_inst[15:11] == 5'b10011 &&
	      fn_decompress_inst[6:0] == 7'b0000010 ||
	      fn_decompress_inst[15:12] == 4'b1001 &&
	      fn_decompress_inst_BIT_10_AND_fn_decompress_in_ETC___d277) ?
	       { 12'd0, fn_decompress_inst[11:7], 15'd231 } :
	       IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1001__ETC___d318 ;
  assign IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d322 =
	     (fn_decompress_inst[15:11] == 5'b10001 &&
	      fn_decompress_inst[6:0] == 7'b0000010 ||
	      fn_decompress_inst[15:12] == 4'b1000 &&
	      fn_decompress_inst_BIT_10_AND_fn_decompress_in_ETC___d277) ?
	       { 12'd0, fn_decompress_inst[11:7], 15'd103 } :
	       IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1000__ETC___d321 ;
  assign IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1000__ETC___d321 =
	     (fn_decompress_inst[15:12] == 4'b1000 &&
	      (fn_decompress_inst[6] && fn_decompress_inst[1:0] == 2'b10 ||
	       fn_decompress_inst_BIT_5_4_AND_fn_decompress_i_ETC___d288)) ?
	       { 7'b0,
		 fn_decompress_inst[6:2],
		 8'd0,
		 fn_decompress_inst[11:7],
		 7'd51 } :
	       ((fn_decompress_inst == 16'b1001000000000010) ?
		  32'd1048691 :
		  IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d319) ;
  assign IF_fn_decompress_inst_BITS_15_TO_12_EQ_0b1001__ETC___d318 =
	     (fn_decompress_inst[15:12] == 4'b1001 &&
	      (fn_decompress_inst[6] && fn_decompress_inst[1:0] == 2'b10 ||
	       fn_decompress_inst_BIT_5_4_AND_fn_decompress_i_ETC___d288)) ?
	       { 7'b0,
		 fn_decompress_inst[6:2],
		 fn_decompress_inst[11:7],
		 3'b0,
		 fn_decompress_inst[11:7],
		 7'd51 } :
	       IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b110_8_ETC___d317 ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b100_8_ETC___d335 =
	     (fn_decompress_inst[15:13] == 3'b100 &&
	      fn_decompress_inst[11:10] == 2'b10 &&
	      fn_decompress_inst[1:0] == 2'b01) ?
	       { SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67,
		 2'b01,
		 fn_decompress_inst[9:7],
		 5'b11101,
		 fn_decompress_inst[9:7],
		 7'd19 } :
	       ((fn_decompress_inst[15:10] == 6'b100011 &&
		 fn_decompress_inst[6:5] == 2'b0 &&
		 fn_decompress_inst[1:0] == 2'b01) ?
		  { 9'b010000001,
		    fn_decompress_inst[4:2],
		    2'b01,
		    fn_decompress_inst[9:7],
		    5'b00001,
		    fn_decompress_inst[9:7],
		    7'd51 } :
		  ((fn_decompress_inst[15:10] == 6'b100011 &&
		    fn_decompress_inst[6:5] == 2'b01 &&
		    fn_decompress_inst[1:0] == 2'b01) ?
		     { 9'b000000001,
		       fn_decompress_inst[4:2],
		       2'b01,
		       fn_decompress_inst[9:7],
		       5'b10001,
		       fn_decompress_inst[9:7],
		       7'd51 } :
		     ((fn_decompress_inst[15:10] == 6'b100011 &&
		       fn_decompress_inst[6:5] == 2'b10 &&
		       fn_decompress_inst[1:0] == 2'b01) ?
			{ 9'b000000001,
			  fn_decompress_inst[4:2],
			  2'b01,
			  fn_decompress_inst[9:7],
			  5'b11001,
			  fn_decompress_inst[9:7],
			  7'd51 } :
			((fn_decompress_inst[15:10] == 6'b100011 &&
			  fn_decompress_inst[6:5] == 2'b11 &&
			  fn_decompress_inst[1:0] == 2'b01) ?
			   { 9'b000000001,
			     fn_decompress_inst[4:2],
			     2'b01,
			     fn_decompress_inst[9:7],
			     5'b11101,
			     fn_decompress_inst[9:7],
			     7'd51 } :
			   ((fn_decompress_inst[15:10] == 6'b100111 &&
			     fn_decompress_inst[6:5] == 2'b0 &&
			     fn_decompress_inst[1:0] == 2'b01) ?
			      { 9'b010000001,
				fn_decompress_inst[4:2],
				2'b01,
				fn_decompress_inst[9:7],
				5'b00001,
				fn_decompress_inst[9:7],
				7'd59 } :
			      ((fn_decompress_inst[15:10] == 6'b100111 &&
				fn_decompress_inst[6:5] == 2'b01 &&
				fn_decompress_inst[1:0] == 2'b01) ?
				 { 9'b000000001,
				   fn_decompress_inst[4:2],
				   2'b01,
				   fn_decompress_inst[9:7],
				   5'b00001,
				   fn_decompress_inst[9:7],
				   7'd59 } :
				 ((fn_decompress_inst[15:13] == 3'b101 &&
				   fn_decompress_inst[1:0] == 2'b01) ?
				    { fn_decompress_inst[12],
				      fn_decompress_inst[8],
				      fn_decompress_inst[10:9],
				      fn_decompress_inst[6],
				      fn_decompress_inst[7],
				      fn_decompress_inst[2],
				      fn_decompress_inst[11],
				      fn_decompress_inst[5:3],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      fn_decompress_inst[12],
				      12'd111 } :
				    ((fn_decompress_inst[15:13] == 3'b110 &&
				      fn_decompress_inst[1:0] == 2'b01) ?
				       { fn_decompress_inst[12],
					 fn_decompress_inst[12],
					 fn_decompress_inst[12],
					 fn_decompress_inst[12],
					 fn_decompress_inst[6:5],
					 fn_decompress_inst[2],
					 7'b0000001,
					 fn_decompress_inst[9:7],
					 3'b0,
					 fn_decompress_inst[11:10],
					 fn_decompress_inst[4:3],
					 fn_decompress_inst[12],
					 7'd99 } :
				       ((fn_decompress_inst[15:13] ==
					 3'b111 &&
					 fn_decompress_inst[1:0] == 2'b01) ?
					  { fn_decompress_inst[12],
					    fn_decompress_inst[12],
					    fn_decompress_inst[12],
					    fn_decompress_inst[12],
					    fn_decompress_inst[6:5],
					    fn_decompress_inst[2],
					    7'b0000001,
					    fn_decompress_inst[9:7],
					    3'b001,
					    fn_decompress_inst[11:10],
					    fn_decompress_inst[4:3],
					    fn_decompress_inst[12],
					    7'd99 } :
					  ((fn_decompress_inst[15:13] ==
					    3'b0 &&
					    fn_decompress_inst[1:0] ==
					    2'b10) ?
					     { 6'b0,
					       fn_decompress_inst[12],
					       fn_decompress_inst[6:2],
					       fn_decompress_inst[11:7],
					       3'b001,
					       fn_decompress_inst[11:7],
					       7'd19 } :
					     IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b10_2__ETC___d324)))))))))) ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b10_2__ETC___d324 =
	     (fn_decompress_inst[15:13] == 3'b010 &&
	      (fn_decompress_inst[11] || fn_decompress_inst[10] ||
	       fn_decompress_inst[9] ||
	       fn_decompress_inst[8] ||
	       fn_decompress_inst[7]) &&
	      fn_decompress_inst[1:0] == 2'b10) ?
	       { 4'd0, x__h12096, 8'd18, fn_decompress_inst[11:7], 7'd3 } :
	       ((fn_decompress_inst[15:13] == 3'b011 &&
		 fn_decompress_inst[1:0] == 2'b10) ?
		  { 3'd0, x__h12235, 8'd19, fn_decompress_inst[11:7], 7'd3 } :
		  IF_fn_decompress_inst_BITS_15_TO_11_11_EQ_0b10_ETC___d322) ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b110_8_ETC___d317 =
	     (fn_decompress_inst[15:13] == 3'b110 &&
	      fn_decompress_inst[1:0] == 2'b10) ?
	       { 4'd0,
		 x__h14479,
		 fn_decompress_inst[6:2],
		 8'd18,
		 fn_decompress_inst[11:9],
		 9'd35 } :
	       ((fn_decompress_inst[15:13] == 3'b111 &&
		 fn_decompress_inst[1:0] == 2'b10) ?
		  { 3'd0,
		    x__h14618,
		    fn_decompress_inst[6:2],
		    8'd19,
		    fn_decompress_inst[11:10],
		    10'd35 } :
		  32'd0) ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b111_7_ETC___d343 =
	     (fn_decompress_inst[15:13] == 3'b111 &&
	      fn_decompress_inst[1:0] == 2'b0) ?
	       { 4'd0,
		 x__h2058,
		 2'b01,
		 fn_decompress_inst[4:2],
		 2'b01,
		 fn_decompress_inst[9:7],
		 3'b011,
		 fn_decompress_inst[11:10],
		 10'd35 } :
	       ((fn_decompress_inst[15:13] == 3'b0 &&
		 fn_decompress_inst[1:0] == 2'b01) ?
		  { SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67,
		    fn_decompress_inst[11:7],
		    3'b0,
		    fn_decompress_inst[11:7],
		    7'd19 } :
		  IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b1_2_A_ETC___d341) ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b11_2__ETC___d345 =
	     (fn_decompress_inst[15:13] == 3'b011 &&
	      fn_decompress_inst[1:0] == 2'b0) ?
	       { 4'd0,
		 x__h1733,
		 2'b01,
		 fn_decompress_inst[9:7],
		 5'b01101,
		 fn_decompress_inst[4:2],
		 7'd3 } :
	       ((fn_decompress_inst[15:13] == 3'b110 &&
		 fn_decompress_inst[1:0] == 2'b0) ?
		  { 5'd0,
		    x__h1873,
		    2'b01,
		    fn_decompress_inst[4:2],
		    2'b01,
		    fn_decompress_inst[9:7],
		    3'b010,
		    fn_decompress_inst[11:10],
		    fn_decompress_inst[6],
		    9'd35 } :
		  IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b111_7_ETC___d343) ;
  assign IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b1_2_A_ETC___d341 =
	     (fn_decompress_inst[15:13] == 3'b001 &&
	      (fn_decompress_inst[11] || fn_decompress_inst[10] ||
	       fn_decompress_inst[9] ||
	       fn_decompress_inst[8] ||
	       fn_decompress_inst[7]) &&
	      fn_decompress_inst[1:0] == 2'b01) ?
	       { SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67,
		 fn_decompress_inst[11:7],
		 3'b0,
		 fn_decompress_inst[11:7],
		 7'd27 } :
	       ((fn_decompress_inst[15:13] == 3'b010 &&
		 fn_decompress_inst[1:0] == 2'b01) ?
		  { SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67,
		    8'd0,
		    fn_decompress_inst[11:7],
		    7'd19 } :
		  IF_fn_decompress_inst_BITS_15_TO_7_3_EQ_0b1110_ETC___d339) ;
  assign IF_fn_decompress_inst_BITS_15_TO_7_3_EQ_0b1110_ETC___d339 =
	     (fn_decompress_inst[15:7] == 9'b011100010 &&
	      fn_decompress_inst[1:0] == 2'b01 ||
	      fn_decompress_inst[15:13] == 3'b011 &&
	      (fn_decompress_inst[11:6] == 6'b000101 &&
	       fn_decompress_inst[1:0] == 2'b01 ||
	       fn_decompress_inst[11:7] == 5'b00010 &&
	       (fn_decompress_inst[5] && fn_decompress_inst[1:0] == 2'b01 ||
		fn_decompress_inst[4] && fn_decompress_inst[1:0] == 2'b01 ||
		fn_decompress_inst[3] && fn_decompress_inst[1:0] == 2'b01 ||
		fn_decompress_inst[2:0] == 3'b101))) ?
	       { { {2{x__h4254[9]}}, x__h4254 }, 20'd65811 } :
	       ((fn_decompress_inst[15:11] == 5'b01111 &&
		 fn_decompress_inst[1:0] == 2'b01 ||
		 fn_decompress_inst[15:12] == 4'b0111 &&
		 fn_decompress_inst[10] &&
		 fn_decompress_inst[1:0] == 2'b01 ||
		 fn_decompress_inst[15:12] == 4'b0111 &&
		 fn_decompress_inst[9] &&
		 fn_decompress_inst[1:0] == 2'b01 ||
		 fn_decompress_inst[15:12] == 4'b0111 &&
		 !fn_decompress_inst[8] &&
		 fn_decompress_inst[1:0] == 2'b01 ||
		 fn_decompress_inst[15:12] == 4'b0111 &&
		 fn_decompress_inst[7] &&
		 fn_decompress_inst[1:0] == 2'b01 ||
		 fn_decompress_inst[15:13] == 3'b011 &&
		 (fn_decompress_inst[11] && fn_decompress_inst[6] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[10] && fn_decompress_inst[6] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[9] && fn_decompress_inst[6] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  !fn_decompress_inst[8] && fn_decompress_inst[6] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[7:6] == 2'b11 &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[11] && fn_decompress_inst[5] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[10] && fn_decompress_inst[5] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[9] && fn_decompress_inst[5] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  !fn_decompress_inst[8] && fn_decompress_inst[5] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[7] && fn_decompress_inst[5] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[11] && fn_decompress_inst[4] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[10] && fn_decompress_inst[4] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[9] && fn_decompress_inst[4] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  !fn_decompress_inst[8] && fn_decompress_inst[4] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[7] && fn_decompress_inst[4] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[11] && fn_decompress_inst[3] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[10] && fn_decompress_inst[3] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[9] && fn_decompress_inst[3] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  !fn_decompress_inst[8] && fn_decompress_inst[3] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  fn_decompress_inst[7] && fn_decompress_inst[3] &&
		  fn_decompress_inst[1:0] == 2'b01 ||
		  (fn_decompress_inst[11] || fn_decompress_inst[10] ||
		   fn_decompress_inst[9] ||
		   !fn_decompress_inst[8] ||
		   fn_decompress_inst[7]) &&
		  fn_decompress_inst[2:0] == 3'b101)) ?
		  { { {14{fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1[5]}},
		      fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1 },
		    fn_decompress_inst[11:7],
		    7'd55 } :
		  ((fn_decompress_inst[15:13] == 3'b100 &&
		    fn_decompress_inst[11:10] == 2'b0 &&
		    fn_decompress_inst[1:0] == 2'b01) ?
		     { 6'b0,
		       fn_decompress_inst[12],
		       fn_decompress_inst[6:2],
		       2'b01,
		       fn_decompress_inst[9:7],
		       5'b10101,
		       fn_decompress_inst[9:7],
		       7'd19 } :
		     ((fn_decompress_inst[15:13] == 3'b100 &&
		       fn_decompress_inst[11:10] == 2'b01 &&
		       fn_decompress_inst[1:0] == 2'b01) ?
			{ 6'b010000,
			  fn_decompress_inst[12],
			  fn_decompress_inst[6:2],
			  2'b01,
			  fn_decompress_inst[9:7],
			  5'b10101,
			  fn_decompress_inst[9:7],
			  7'd19 } :
			IF_fn_decompress_inst_BITS_15_TO_13_EQ_0b100_8_ETC___d335))) ;
  assign SEXT_fn_decompress_inst_BIT_12_0_CONCAT_fn_dec_ETC___d67 =
	     { {6{fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1[5]}},
	       fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1 } ;
  assign fn_decompress_inst_BIT_10_AND_fn_decompress_in_ETC___d277 =
	     fn_decompress_inst[10] &&
	     fn_decompress_inst[6:0] == 7'b0000010 ||
	     fn_decompress_inst[9] && fn_decompress_inst[6:0] == 7'b0000010 ||
	     fn_decompress_inst[8] && fn_decompress_inst[6:0] == 7'b0000010 ||
	     fn_decompress_inst[7:0] == 8'b10000010 ;
  assign fn_decompress_inst_BIT_12_CONCAT_fn_decompress_ETC__q1 =
	     { fn_decompress_inst[12], fn_decompress_inst[6:2] } ;
  assign fn_decompress_inst_BIT_5_4_AND_fn_decompress_i_ETC___d288 =
	     fn_decompress_inst[5] && fn_decompress_inst[1:0] == 2'b10 ||
	     fn_decompress_inst[4] && fn_decompress_inst[1:0] == 2'b10 ||
	     fn_decompress_inst[3] && fn_decompress_inst[1:0] == 2'b10 ||
	     fn_decompress_inst[2:0] == 3'b110 ;
  assign x__h12096 =
	     { fn_decompress_inst[3:2],
	       fn_decompress_inst[12],
	       fn_decompress_inst[6:4],
	       2'd0 } ;
  assign x__h12235 =
	     { fn_decompress_inst[4:2],
	       fn_decompress_inst[12],
	       fn_decompress_inst[6:5],
	       3'd0 } ;
  assign x__h1408 =
	     { fn_decompress_inst[10:7],
	       fn_decompress_inst[12:11],
	       fn_decompress_inst[5],
	       fn_decompress_inst[6],
	       2'd0 } ;
  assign x__h14479 = { fn_decompress_inst[8:7], fn_decompress_inst[12] } ;
  assign x__h14618 = { fn_decompress_inst[9:7], fn_decompress_inst[12] } ;
  assign x__h1569 =
	     { fn_decompress_inst[5],
	       fn_decompress_inst[12:10],
	       fn_decompress_inst[6],
	       2'd0 } ;
  assign x__h1733 =
	     { fn_decompress_inst[6:5], fn_decompress_inst[12:10], 3'd0 } ;
  assign x__h1873 = { fn_decompress_inst[5], fn_decompress_inst[12] } ;
  assign x__h2058 = { fn_decompress_inst[6:5], fn_decompress_inst[12] } ;
  assign x__h4254 =
	     { fn_decompress_inst[12],
	       fn_decompress_inst[4:3],
	       fn_decompress_inst[5],
	       fn_decompress_inst[2],
	       fn_decompress_inst[6],
	       4'd0 } ;
endmodule  // module_fn_decompress

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:36:51 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// fn_pmp_lookup                  O     7
// fn_pmp_lookup_req              I    40
// fn_pmp_lookup_priv             I     2
// fn_pmp_lookup_pmpcfg           I    32
// fn_pmp_lookup_pmpaddr          I   120
//
// Combinational paths from inputs to outputs:
//   (fn_pmp_lookup_req,
//    fn_pmp_lookup_priv,
//    fn_pmp_lookup_pmpcfg,
//    fn_pmp_lookup_pmpaddr) -> fn_pmp_lookup
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_fn_pmp_lookup(fn_pmp_lookup_req,
			    fn_pmp_lookup_priv,
			    fn_pmp_lookup_pmpcfg,
			    fn_pmp_lookup_pmpaddr,
			    fn_pmp_lookup);
  // value method fn_pmp_lookup
  input  [39 : 0] fn_pmp_lookup_req;
  input  [1 : 0] fn_pmp_lookup_priv;
  input  [31 : 0] fn_pmp_lookup_pmpcfg;
  input  [119 : 0] fn_pmp_lookup_pmpaddr;
  output [6 : 0] fn_pmp_lookup;

  // signals for module outputs
  wire [6 : 0] fn_pmp_lookup;

  // remaining internal signals
  reg [5 : 0] x__h10555;
  reg IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168,
      IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361,
      IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252,
      IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375,
      IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336,
      IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348,
      IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85;
  wire [31 : 0] mask__h3039,
		mask__h437,
		mask__h5349,
		mask__h7659,
		reqtop__h30,
		x__h3121,
		x__h3207,
		x__h5431,
		x__h5517,
		x__h7741,
		x__h7827,
		x__h897,
		y__h2991,
		y__h3208,
		y__h5300,
		y__h5518,
		y__h7610,
		y__h7770,
		y__h7828,
		y__h898,
		y__h9920;
  wire [29 : 0] INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4,
		INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1,
		INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2,
		INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3;
  wire [4 : 0] x__h2986, x__h5295, x__h7605, x__h9915;
  wire IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d378,
       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d379,
       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d444,
       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d445,
       fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11,
       fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79,
       fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81,
       fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88,
       fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162,
       fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164,
       fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172,
       fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94,
       fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178,
       fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246,
       fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91,
       fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95;

  // value method fn_pmp_lookup
  assign fn_pmp_lookup =
	     { (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85 ||
		IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168 ||
		IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252 ||
		IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336) &&
	       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d379 &&
	       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d445,
	       x__h10555 } ;

  // remaining internal signals
  assign IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d378 =
	     (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361) ?
	       IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252 :
	       (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 ?
		  IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168 :
		  IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85) ;
  assign IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d379 =
	     (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375) ?
	       IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336 :
	       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d378 ;
  assign IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d444 =
	     (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361) ?
	       (fn_pmp_lookup_pmpcfg[23] || fn_pmp_lookup_priv != 2'd3) &&
	       (fn_pmp_lookup_req[1:0] == 2'd0 && !fn_pmp_lookup_pmpcfg[16] ||
		fn_pmp_lookup_req[1:0] == 2'd1 && !fn_pmp_lookup_pmpcfg[17] ||
		fn_pmp_lookup_req[1:0] == 2'd2 && !fn_pmp_lookup_pmpcfg[18]) :
	       (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 ?
		  (fn_pmp_lookup_pmpcfg[15] || fn_pmp_lookup_priv != 2'd3) &&
		  (fn_pmp_lookup_req[1:0] == 2'd0 &&
		   !fn_pmp_lookup_pmpcfg[8] ||
		   fn_pmp_lookup_req[1:0] == 2'd1 &&
		   !fn_pmp_lookup_pmpcfg[9] ||
		   fn_pmp_lookup_req[1:0] == 2'd2 &&
		   !fn_pmp_lookup_pmpcfg[10]) :
		  (fn_pmp_lookup_pmpcfg[7] || fn_pmp_lookup_priv != 2'd3) &&
		  (fn_pmp_lookup_req[1:0] == 2'd0 &&
		   !fn_pmp_lookup_pmpcfg[0] ||
		   fn_pmp_lookup_req[1:0] == 2'd1 &&
		   !fn_pmp_lookup_pmpcfg[1] ||
		   fn_pmp_lookup_req[1:0] == 2'd2 &&
		   !fn_pmp_lookup_pmpcfg[2])) ;
  assign IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d445 =
	     (IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361 &&
	      IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375) ?
	       (fn_pmp_lookup_pmpcfg[31] || fn_pmp_lookup_priv != 2'd3) &&
	       (fn_pmp_lookup_req[1:0] == 2'd0 && !fn_pmp_lookup_pmpcfg[24] ||
		fn_pmp_lookup_req[1:0] == 2'd1 && !fn_pmp_lookup_pmpcfg[25] ||
		fn_pmp_lookup_req[1:0] == 2'd2 && !fn_pmp_lookup_pmpcfg[26]) :
	       IF_IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_TH_ETC___d444 ;
  assign INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4 =
	     ~fn_pmp_lookup_pmpaddr[119:90] ;
  assign INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1 =
	     ~fn_pmp_lookup_pmpaddr[29:0] ;
  assign INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2 =
	     ~fn_pmp_lookup_pmpaddr[59:30] ;
  assign INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3 =
	     ~fn_pmp_lookup_pmpaddr[89:60] ;
  assign fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11 =
	     x__h3121 == fn_pmp_lookup_req[39:8] ;
  assign fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79 =
	     x__h897 == y__h898 ;
  assign fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81 =
	     x__h897 == y__h2991 ;
  assign fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88 =
	     x__h3121 <= fn_pmp_lookup_req[39:8] ;
  assign fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162 =
	     x__h3207 == y__h3208 ;
  assign fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164 =
	     x__h3207 == y__h5300 ;
  assign fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172 =
	     x__h5431 <= fn_pmp_lookup_req[39:8] ;
  assign fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94 =
	     x__h5431 == fn_pmp_lookup_req[39:8] ;
  assign fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178 =
	     x__h7741 == fn_pmp_lookup_req[39:8] ;
  assign fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246 =
	     x__h5517 == y__h5518 ;
  assign fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248 =
	     x__h5517 == y__h7610 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12 =
	     reqtop__h30 == x__h3121 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175 =
	     reqtop__h30 <= x__h7741 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179 =
	     reqtop__h30 == x__h7741 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9 =
	     reqtop__h30 <= x__h3121 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91 =
	     reqtop__h30 <= x__h5431 ;
  assign fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95 =
	     reqtop__h30 == x__h5431 ;
  assign mask__h3039 = 32'hFFFFFFF8 << x__h5295 ;
  assign mask__h437 = 32'hFFFFFFF8 << x__h2986 ;
  assign mask__h5349 = 32'hFFFFFFF8 << x__h7605 ;
  assign mask__h7659 = 32'hFFFFFFF8 << x__h9915 ;
  assign reqtop__h30 =
	     fn_pmp_lookup_req[39:8] + { 26'd0, fn_pmp_lookup_req[7:2] } ;
  assign x__h2986 =
	     INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[0] ?
	       5'd0 :
	       (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[1] ?
		  5'd1 :
		  (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[2] ?
		     5'd2 :
		     (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[3] ?
			5'd3 :
			(INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[4] ?
			   5'd4 :
			   (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[5] ?
			      5'd5 :
			      (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[6] ?
				 5'd6 :
				 (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[7] ?
				    5'd7 :
				    (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[8] ?
				       5'd8 :
				       (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[9] ?
					  5'd9 :
					  (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[10] ?
					     5'd10 :
					     (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[11] ?
						5'd11 :
						(INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[12] ?
						   5'd12 :
						   (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[13] ?
						      5'd13 :
						      (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[14] ?
							 5'd14 :
							 (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[15] ?
							    5'd15 :
							    (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[16] ?
							       5'd16 :
							       (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[17] ?
								  5'd17 :
								  (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[18] ?
								     5'd18 :
								     (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[19] ?
									5'd19 :
									(INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[20] ?
									   5'd20 :
									   (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[21] ?
									      5'd21 :
									      (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[22] ?
										 5'd22 :
										 (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[23] ?
										    5'd23 :
										    (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[24] ?
										       5'd24 :
										       (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[25] ?
											  5'd25 :
											  (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[26] ?
											     5'd26 :
											     (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[27] ?
												5'd27 :
												(INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[28] ?
												   5'd28 :
												   (INV_fn_pmp_lookup_pmpaddr_BITS_29_TO_0__q1[29] ?
												      5'd29 :
												      5'd30))))))))))))))))))))))))))))) ;
  assign x__h3121 = { fn_pmp_lookup_pmpaddr[29:0], 2'b0 } ;
  assign x__h3207 = x__h5431 & mask__h3039 ;
  assign x__h5295 =
	     INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[0] ?
	       5'd0 :
	       (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[1] ?
		  5'd1 :
		  (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[2] ?
		     5'd2 :
		     (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[3] ?
			5'd3 :
			(INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[4] ?
			   5'd4 :
			   (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[5] ?
			      5'd5 :
			      (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[6] ?
				 5'd6 :
				 (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[7] ?
				    5'd7 :
				    (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[8] ?
				       5'd8 :
				       (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[9] ?
					  5'd9 :
					  (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[10] ?
					     5'd10 :
					     (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[11] ?
						5'd11 :
						(INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[12] ?
						   5'd12 :
						   (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[13] ?
						      5'd13 :
						      (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[14] ?
							 5'd14 :
							 (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[15] ?
							    5'd15 :
							    (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[16] ?
							       5'd16 :
							       (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[17] ?
								  5'd17 :
								  (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[18] ?
								     5'd18 :
								     (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[19] ?
									5'd19 :
									(INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[20] ?
									   5'd20 :
									   (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[21] ?
									      5'd21 :
									      (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[22] ?
										 5'd22 :
										 (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[23] ?
										    5'd23 :
										    (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[24] ?
										       5'd24 :
										       (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[25] ?
											  5'd25 :
											  (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[26] ?
											     5'd26 :
											     (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[27] ?
												5'd27 :
												(INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[28] ?
												   5'd28 :
												   (INV_fn_pmp_lookup_pmpaddr_BITS_59_TO_30__q2[29] ?
												      5'd29 :
												      5'd30))))))))))))))))))))))))))))) ;
  assign x__h5431 = { fn_pmp_lookup_pmpaddr[59:30], 2'b0 } ;
  assign x__h5517 = x__h7741 & mask__h5349 ;
  assign x__h7605 =
	     INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[0] ?
	       5'd0 :
	       (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[1] ?
		  5'd1 :
		  (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[2] ?
		     5'd2 :
		     (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[3] ?
			5'd3 :
			(INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[4] ?
			   5'd4 :
			   (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[5] ?
			      5'd5 :
			      (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[6] ?
				 5'd6 :
				 (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[7] ?
				    5'd7 :
				    (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[8] ?
				       5'd8 :
				       (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[9] ?
					  5'd9 :
					  (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[10] ?
					     5'd10 :
					     (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[11] ?
						5'd11 :
						(INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[12] ?
						   5'd12 :
						   (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[13] ?
						      5'd13 :
						      (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[14] ?
							 5'd14 :
							 (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[15] ?
							    5'd15 :
							    (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[16] ?
							       5'd16 :
							       (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[17] ?
								  5'd17 :
								  (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[18] ?
								     5'd18 :
								     (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[19] ?
									5'd19 :
									(INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[20] ?
									   5'd20 :
									   (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[21] ?
									      5'd21 :
									      (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[22] ?
										 5'd22 :
										 (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[23] ?
										    5'd23 :
										    (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[24] ?
										       5'd24 :
										       (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[25] ?
											  5'd25 :
											  (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[26] ?
											     5'd26 :
											     (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[27] ?
												5'd27 :
												(INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[28] ?
												   5'd28 :
												   (INV_fn_pmp_lookup_pmpaddr_BITS_89_TO_60__q3[29] ?
												      5'd29 :
												      5'd30))))))))))))))))))))))))))))) ;
  assign x__h7741 = { fn_pmp_lookup_pmpaddr[89:60], 2'b0 } ;
  assign x__h7827 = y__h7770 & mask__h7659 ;
  assign x__h897 = x__h3121 & mask__h437 ;
  assign x__h9915 =
	     INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[0] ?
	       5'd0 :
	       (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[1] ?
		  5'd1 :
		  (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[2] ?
		     5'd2 :
		     (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[3] ?
			5'd3 :
			(INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[4] ?
			   5'd4 :
			   (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[5] ?
			      5'd5 :
			      (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[6] ?
				 5'd6 :
				 (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[7] ?
				    5'd7 :
				    (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[8] ?
				       5'd8 :
				       (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[9] ?
					  5'd9 :
					  (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[10] ?
					     5'd10 :
					     (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[11] ?
						5'd11 :
						(INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[12] ?
						   5'd12 :
						   (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[13] ?
						      5'd13 :
						      (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[14] ?
							 5'd14 :
							 (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[15] ?
							    5'd15 :
							    (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[16] ?
							       5'd16 :
							       (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[17] ?
								  5'd17 :
								  (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[18] ?
								     5'd18 :
								     (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[19] ?
									5'd19 :
									(INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[20] ?
									   5'd20 :
									   (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[21] ?
									      5'd21 :
									      (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[22] ?
										 5'd22 :
										 (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[23] ?
										    5'd23 :
										    (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[24] ?
										       5'd24 :
										       (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[25] ?
											  5'd25 :
											  (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[26] ?
											     5'd26 :
											     (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[27] ?
												5'd27 :
												(INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[28] ?
												   5'd28 :
												   (INV_fn_pmp_lookup_pmpaddr_BITS_119_TO_90__q4[29] ?
												      5'd29 :
												      5'd30))))))))))))))))))))))))))))) ;
  assign y__h2991 = reqtop__h30 & mask__h437 ;
  assign y__h3208 = fn_pmp_lookup_req[39:8] & mask__h3039 ;
  assign y__h5300 = reqtop__h30 & mask__h3039 ;
  assign y__h5518 = fn_pmp_lookup_req[39:8] & mask__h5349 ;
  assign y__h7610 = reqtop__h30 & mask__h5349 ;
  assign y__h7770 = { fn_pmp_lookup_pmpaddr[119:90], 2'b0 } ;
  assign y__h7828 = fn_pmp_lookup_req[39:8] & mask__h7659 ;
  assign y__h898 = fn_pmp_lookup_req[39:8] & mask__h437 ;
  assign y__h9920 = reqtop__h30 & mask__h7659 ;
  always@(fn_pmp_lookup_req)
  begin
    case (fn_pmp_lookup_req[1:0])
      2'd0: x__h10555 = 6'd5;
      2'd1: x__h10555 = 6'd7;
      default: x__h10555 = 6'd1;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12)
  begin
    case (fn_pmp_lookup_pmpcfg[4:3])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85 =
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85 =
	      fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11 &&
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d85 =
		   fn_pmp_lookup_pmpcfg[4:3] == 2'd3 &&
		   fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79 &&
		   fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95)
  begin
    case (fn_pmp_lookup_pmpcfg[12:11])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168 =
	      fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88 &&
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168 =
	      fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94 &&
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d168 =
		   fn_pmp_lookup_pmpcfg[12:11] == 2'd3 &&
		   fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162 &&
		   fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246 or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175 or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179)
  begin
    case (fn_pmp_lookup_pmpcfg[20:19])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252 =
	      fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172 &&
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252 =
	      fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178 &&
	      fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d252 =
		   fn_pmp_lookup_pmpcfg[20:19] == 2'd3 &&
		   fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246 &&
		   fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12)
  begin
    case (fn_pmp_lookup_pmpcfg[4:3])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 =
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d9;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 =
	      !fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d11 ||
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d12;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_4_TO_3_EQ_1_THEN__ETC___d348 =
		   fn_pmp_lookup_pmpcfg[4:3] != 2'd3 ||
		   !fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d79 ||
		   !fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d81;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164 or
	  fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95)
  begin
    case (fn_pmp_lookup_pmpcfg[12:11])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361 =
	      !fn_pmp_lookup_pmpaddr_BITS_29_TO_0_CONCAT_0b0__ETC___d88 ||
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d91;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361 =
	      !fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d94 ||
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d95;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_12_TO_11_6_EQ_1_7_ETC___d361 =
		   fn_pmp_lookup_pmpcfg[12:11] != 2'd3 ||
		   !fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d162 ||
		   !fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d164;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246 or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248 or
	  fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175 or
	  fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178 or
	  fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179)
  begin
    case (fn_pmp_lookup_pmpcfg[20:19])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375 =
	      !fn_pmp_lookup_pmpaddr_BITS_59_TO_30_9_CONCAT_0_ETC___d172 ||
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d175;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375 =
	      !fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d178 ||
	      !fn_pmp_lookup_req_BITS_39_TO_8_PLUS_0_CONCAT_f_ETC___d179;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_20_TO_19_70_EQ_1__ETC___d375 =
		   fn_pmp_lookup_pmpcfg[20:19] != 2'd3 ||
		   !fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d246 ||
		   !fn_pmp_lookup_pmpaddr_BITS_89_TO_60_73_CONCAT__ETC___d248;
    endcase
  end
  always@(fn_pmp_lookup_pmpcfg or
	  x__h7827 or
	  y__h7828 or
	  y__h9920 or
	  x__h7741 or fn_pmp_lookup_req or reqtop__h30 or y__h7770)
  begin
    case (fn_pmp_lookup_pmpcfg[28:27])
      2'd1:
	  IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336 =
	      x__h7741 <= fn_pmp_lookup_req[39:8] && reqtop__h30 <= y__h7770;
      2'd2:
	  IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336 =
	      y__h7770 == fn_pmp_lookup_req[39:8] && reqtop__h30 == y__h7770;
      default: IF_fn_pmp_lookup_pmpcfg_BITS_28_TO_27_54_EQ_1__ETC___d336 =
		   fn_pmp_lookup_pmpcfg[28:27] == 2'd3 &&
		   x__h7827 == y__h7828 &&
		   x__h7827 == y__h9920;
    endcase
  end
endmodule  // module_fn_pmp_lookup

//
// Generated by Bluespec Compiler, version 2018.10.beta1 (build e1df8052c, 2018-10-17)
//
// On Tue Oct  1 16:37:12 IST 2019
//
//
// Ports:
// Name                         I/O  size props
// singlestep                     O   129
// singlestep_remainder           I    65
// singlestep_quotient            I    64
// singlestep_divisor             I    64
//
// Combinational paths from inputs to outputs:
//   (singlestep_remainder,
//    singlestep_quotient,
//    singlestep_divisor) -> singlestep
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module module_singlestep(singlestep_remainder,
			 singlestep_quotient,
			 singlestep_divisor,
			 singlestep);
  // value method singlestep
  input  [64 : 0] singlestep_remainder;
  input  [63 : 0] singlestep_quotient;
  input  [63 : 0] singlestep_divisor;
  output [128 : 0] singlestep;

  // signals for module outputs
  wire [128 : 0] singlestep;

  // remaining internal signals
  wire [64 : 0] remainder__h62, sub__h64, x__h24;
  wire [63 : 0] x__h101, x__h96;
  wire singlestep_remainder_BITS_62_TO_0_CONCAT_singl_ETC___d4;

  // value method singlestep
  assign singlestep = { x__h24, x__h101 } ;

  // remaining internal signals
  assign remainder__h62 =
	     { singlestep_remainder[63:0], singlestep_quotient[63] } ;
  assign singlestep_remainder_BITS_62_TO_0_CONCAT_singl_ETC___d4 =
	     { singlestep_remainder[62:0], singlestep_quotient[63] } <
	     singlestep_divisor ;
  assign sub__h64 = remainder__h62 + { x__h96[63], x__h96 } ;
  assign x__h101 =
	     { singlestep_quotient[62:0],
	       !singlestep_remainder_BITS_62_TO_0_CONCAT_singl_ETC___d4 } ;
  assign x__h24 =
	     singlestep_remainder_BITS_62_TO_0_CONCAT_singl_ETC___d4 ?
	       remainder__h62 :
	       sub__h64 ;
  assign x__h96 = ~singlestep_divisor + 64'd1 ;
endmodule  // module_singlestep


// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision: 24080 $
// $Date: 2011-05-18 15:32:52 -0400 (Wed, 18 May 2011) $

`ifdef  BSV_WARN_REGFILE_ADDR_RANGE
`else
`define BSV_WARN_REGFILE_ADDR_RANGE 0
`endif

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif


// Multi-ported Register File -- initializable from a file.
module RegFileLoad(CLK,
                   ADDR_IN, D_IN, WE,
                   ADDR_1, D_OUT_1,
                   ADDR_2, D_OUT_2,
                   ADDR_3, D_OUT_3,
                   ADDR_4, D_OUT_4,
                   ADDR_5, D_OUT_5
                   );
   parameter                   file = "";
   parameter                   addr_width = 1;
   parameter                   data_width = 1;
   parameter                   lo = 0;
   parameter                   hi = 1;
   parameter                   binary = 0;

   input                       CLK;
   input [addr_width - 1 : 0]  ADDR_IN;
   input [data_width - 1 : 0]  D_IN;
   input                       WE;

   input [addr_width - 1 : 0]  ADDR_1;
   output [data_width - 1 : 0] D_OUT_1;

   input [addr_width - 1 : 0]  ADDR_2;
   output [data_width - 1 : 0] D_OUT_2;

   input [addr_width - 1 : 0]  ADDR_3;
   output [data_width - 1 : 0] D_OUT_3;

   input [addr_width - 1 : 0]  ADDR_4;
   output [data_width - 1 : 0] D_OUT_4;

   input [addr_width - 1 : 0]  ADDR_5;
   output [data_width - 1 : 0] D_OUT_5;

   reg [data_width - 1 : 0]    arr[lo:hi];


   initial
     begin : init_rom_block
	if (binary)
           $readmemb(file, arr, lo, hi);
        else
           $readmemh(file, arr, lo, hi);
     end // initial begin


   always@(posedge CLK)
     begin
        if (WE)
          arr[ADDR_IN] <= `BSV_ASSIGNMENT_DELAY D_IN;
     end // always@ (posedge CLK)

   assign D_OUT_1 = arr[ADDR_1];
   assign D_OUT_2 = arr[ADDR_2];
   assign D_OUT_3 = arr[ADDR_3];
   assign D_OUT_4 = arr[ADDR_4];
   assign D_OUT_5 = arr[ADDR_5];

   // synopsys translate_off
   always@(posedge CLK)
     begin : runtime_check
        reg enable_check;
        enable_check = `BSV_WARN_REGFILE_ADDR_RANGE ;
        if ( enable_check )
           begin
              if (( ADDR_1 < lo ) || (ADDR_1 > hi) )
                $display( "Warning: RegFile: %m -- Address port 1 is out of bounds: %h", ADDR_1 ) ;
              if (( ADDR_2 < lo ) || (ADDR_2 > hi) )
                $display( "Warning: RegFile: %m -- Address port 2 is out of bounds: %h", ADDR_2 ) ;
              if (( ADDR_3 < lo ) || (ADDR_3 > hi) )
                $display( "Warning: RegFile: %m -- Address port 3 is out of bounds: %h", ADDR_3 ) ;
              if (( ADDR_4 < lo ) || (ADDR_4 > hi) )
                $display( "Warning: RegFile: %m -- Address port 4 is out of bounds: %h", ADDR_4 ) ;
              if (( ADDR_5 < lo ) || (ADDR_5 > hi) )
                $display( "Warning: RegFile: %m -- Address port 5 is out of bounds: %h", ADDR_5 ) ;
              if ( WE && ( ADDR_IN < lo ) || (ADDR_IN > hi) )
                $display( "Warning: RegFile: %m -- Write Address port is out of bounds: %h", ADDR_IN ) ;
           end
     end
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision: 24080 $
// $Date: 2011-05-18 15:32:52 -0400 (Wed, 18 May 2011) $

`ifdef  BSV_WARN_REGFILE_ADDR_RANGE
`else
`define BSV_WARN_REGFILE_ADDR_RANGE 0 
`endif


`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif


// Multi-ported Register File
module RegFile(CLK,
               ADDR_IN, D_IN, WE,
               ADDR_1, D_OUT_1,
               ADDR_2, D_OUT_2,
               ADDR_3, D_OUT_3,
               ADDR_4, D_OUT_4,
               ADDR_5, D_OUT_5
               );
   parameter                   addr_width = 1;
   parameter                   data_width = 1;
   parameter                   lo = 0;
   parameter                   hi = 1;

   input                       CLK;
   input [addr_width - 1 : 0]  ADDR_IN;
   input [data_width - 1 : 0]  D_IN;
   input                       WE;

   input [addr_width - 1 : 0]  ADDR_1;
   output [data_width - 1 : 0] D_OUT_1;

   input [addr_width - 1 : 0]  ADDR_2;
   output [data_width - 1 : 0] D_OUT_2;

   input [addr_width - 1 : 0]  ADDR_3;
   output [data_width - 1 : 0] D_OUT_3;

   input [addr_width - 1 : 0]  ADDR_4;
   output [data_width - 1 : 0] D_OUT_4;

   input [addr_width - 1 : 0]  ADDR_5;
   output [data_width - 1 : 0] D_OUT_5;

   (* RAM_STYLE = "DISTRIBUTED" *)
   reg [data_width - 1 : 0]    arr[lo:hi];


`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin : init_block
        integer                     i;          // temporary for generate reset value
        for (i = lo; i <= hi; i = i + 1) begin
           arr[i] = {((data_width + 1)/2){2'b10}} ;
        end
     end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


   always@(posedge CLK)
     begin
        if (WE)
          arr[ADDR_IN] <= `BSV_ASSIGNMENT_DELAY D_IN;
     end // always@ (posedge CLK)

   assign D_OUT_1 = arr[ADDR_1];
   assign D_OUT_2 = arr[ADDR_2];
   assign D_OUT_3 = arr[ADDR_3];
   assign D_OUT_4 = arr[ADDR_4];
   assign D_OUT_5 = arr[ADDR_5];

   // synopsys translate_off
   always@(posedge CLK)
     begin : runtime_check
        reg enable_check;
        enable_check = `BSV_WARN_REGFILE_ADDR_RANGE ;
        if ( enable_check )
           begin
              if (( ADDR_1 < lo ) || (ADDR_1 > hi) )
                $display( "Warning: RegFile: %m -- Address port 1 is out of bounds: %h", ADDR_1 ) ;
              if (( ADDR_2 < lo ) || (ADDR_2 > hi) )
                $display( "Warning: RegFile: %m -- Address port 2 is out of bounds: %h", ADDR_2 ) ;
              if (( ADDR_3 < lo ) || (ADDR_3 > hi) )
                $display( "Warning: RegFile: %m -- Address port 3 is out of bounds: %h", ADDR_3 ) ;
              if (( ADDR_4 < lo ) || (ADDR_4 > hi) )
                $display( "Warning: RegFile: %m -- Address port 4 is out of bounds: %h", ADDR_4 ) ;
              if (( ADDR_5 < lo ) || (ADDR_5 > hi) )
                $display( "Warning: RegFile: %m -- Address port 5 is out of bounds: %h", ADDR_5 ) ;
              if ( WE && ( ADDR_IN < lo ) || (ADDR_IN > hi) )
                $display( "Warning: RegFile: %m -- Write Address port is out of bounds: %h", ADDR_IN ) ;
           end
     end
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif



// A separate module which instantiates a simple reset combining primitive.
// The primitive is simply an AND gate for negative resets,  an OR gate for positive resets.
module ResetEither(A_RST,
                   B_RST,
                   RST_OUT
                  ) ;

   input            A_RST;
   input            B_RST;

   output           RST_OUT;

   assign RST_OUT = ((A_RST == `BSV_RESET_VALUE) || (B_RST == `BSV_RESET_VALUE)) ? `BSV_RESET_VALUE : ~ `BSV_RESET_VALUE;

endmodule

// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif

module RevertReg(CLK, Q_OUT, D_IN, EN);

   parameter width = 1;
   parameter init  = { width {1'b0} } ;

   input     CLK;
   input     EN;
   input [width - 1 : 0] D_IN;
   output [width - 1 : 0] Q_OUT;

   assign Q_OUT = init;
endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_ARESET_EDGE_HEAD `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_HEAD
`endif

`ifdef BSV_RESET_FIFO_ARRAY
 `define BSV_ARESET_EDGE_ARRAY `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_ARRAY
`endif


// Sized fifo.  Model has output register which improves timing
module SizedFIFO(CLK, RST, D_IN, ENQ, FULL_N, D_OUT, DEQ, EMPTY_N, CLR);
   parameter               p1width = 1; // data width
   parameter               p2depth = 3;
   parameter               p3cntr_width = 1; // log(p2depth-1)
   // The -1 is allowed since this model has a fast output register
   parameter               guarded = 1;
   localparam              p2depth2 = (p2depth >= 2) ? (p2depth -2) : 0 ;

   input                   CLK;
   input                   RST;
   input                   CLR;
   input [p1width - 1 : 0] D_IN;
   input                   ENQ;
   input                   DEQ;

   output                  FULL_N;
   output                  EMPTY_N;
   output [p1width - 1 : 0] D_OUT;

   reg                      not_ring_full;
   reg                      ring_empty;

   reg [p3cntr_width-1 : 0] head;
   wire [p3cntr_width-1 : 0] next_head;

   reg [p3cntr_width-1 : 0]  tail;
   wire [p3cntr_width-1 : 0] next_tail;

   // if the depth is too small, don't create an ill-sized array;
   // instead, make a 1-sized array and let the initial block report an error
   reg [p1width - 1 : 0]     arr[0: p2depth2];

   reg [p1width - 1 : 0]     D_OUT;
   reg                       hasodata;

   wire [p3cntr_width-1:0]   depthLess2 = p2depth2[p3cntr_width-1:0] ;

   wire [p3cntr_width-1 : 0] incr_tail;
   wire [p3cntr_width-1 : 0] incr_head;

   assign                    incr_tail = tail + 1'b1 ;
   assign                    incr_head = head + 1'b1 ;

   assign    next_head = (head == depthLess2 ) ? {p3cntr_width{1'b0}} : incr_head ;
   assign    next_tail = (tail == depthLess2 ) ? {p3cntr_width{1'b0}} : incr_tail ;

   assign    EMPTY_N = hasodata;
   assign    FULL_N  = not_ring_full;

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin : initial_block
        integer   i;
        D_OUT         = {((p1width + 1)/2){2'b10}} ;

        ring_empty    = 1'b1;
        not_ring_full = 1'b1;
        hasodata      = 1'b0;
        head          = {p3cntr_width {1'b0}} ;
        tail          = {p3cntr_width {1'b0}} ;

        for (i = 0; i <= p2depth2; i = i + 1)
          begin
             arr[i]   = D_OUT ;
          end
     end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


   always @(posedge CLK `BSV_ARESET_EDGE_META)
     begin
        if (RST == `BSV_RESET_VALUE)
          begin
             head <= `BSV_ASSIGNMENT_DELAY {p3cntr_width {1'b0}} ;
             tail <= `BSV_ASSIGNMENT_DELAY {p3cntr_width {1'b0}} ;
             ring_empty <= `BSV_ASSIGNMENT_DELAY 1'b1;
             not_ring_full <= `BSV_ASSIGNMENT_DELAY 1'b1;
             hasodata <= `BSV_ASSIGNMENT_DELAY 1'b0;
          end // if (RST == `BSV_RESET_VALUE)
        else
         begin

             casez ({CLR, DEQ, ENQ, hasodata, ring_empty})
               // Clear operation
               5'b1????: begin
                  head          <= `BSV_ASSIGNMENT_DELAY {p3cntr_width {1'b0}} ;
                  tail          <= `BSV_ASSIGNMENT_DELAY {p3cntr_width {1'b0}} ;
                  ring_empty    <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  not_ring_full <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  hasodata      <= `BSV_ASSIGNMENT_DELAY 1'b0;
               end
               // -----------------------
               // DEQ && ENQ case -- change head and tail if added to ring
               5'b011?0: begin
                  tail          <= `BSV_ASSIGNMENT_DELAY next_tail;
                  head          <= `BSV_ASSIGNMENT_DELAY next_head;
               end
               // -----------------------
               // DEQ only and NO data is in ring
               5'b010?1: begin
                  hasodata <= `BSV_ASSIGNMENT_DELAY 1'b0;
               end
               // DEQ only and data is in ring (move the head pointer)
               5'b010?0: begin
                  head          <= `BSV_ASSIGNMENT_DELAY next_head;
                  not_ring_full <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  ring_empty    <= `BSV_ASSIGNMENT_DELAY next_head == tail ;
               end
               // -----------------------
               // ENQ only when empty
               5'b0010?: begin
                  hasodata      <= `BSV_ASSIGNMENT_DELAY 1'b1;
                  end
               // ENQ only when not empty
               5'b0011?: begin
                  if ( not_ring_full ) // Drop this test to save redundant test
                    // but be warnned that with test fifo overflow causes loss of new data
                    // while without test fifo drops all but head entry! (pointer overflow)
                   begin
                      tail          <= `BSV_ASSIGNMENT_DELAY next_tail;
                      ring_empty    <= `BSV_ASSIGNMENT_DELAY 1'b0;
                      not_ring_full <= `BSV_ASSIGNMENT_DELAY ! (next_tail == head) ;
                   end
               end
             endcase
         end // else: !if(RST == `BSV_RESET_VALUE)
     end // always @ (posedge CLK)

   // Update the fast data out register
   always @(posedge CLK `BSV_ARESET_EDGE_HEAD)
     begin
`ifdef  BSV_RESET_FIFO_HEAD
        if (RST == `BSV_RESET_VALUE)
          begin
             D_OUT    <= `BSV_ASSIGNMENT_DELAY {p1width {1'b0}} ;
          end // if (RST == `BSV_RESET_VALUE)
        else
`endif
        begin
             casez ({CLR, DEQ, ENQ, hasodata, ring_empty})
               // DEQ && ENQ cases
               5'b011?0: begin D_OUT <= `BSV_ASSIGNMENT_DELAY arr[head]; end
               5'b011?1: begin D_OUT <= `BSV_ASSIGNMENT_DELAY D_IN; end
               // DEQ only and data is in ring
               5'b010?0: begin D_OUT <= `BSV_ASSIGNMENT_DELAY arr[head]; end
               // ENQ only when empty
               5'b0010?: begin D_OUT <= `BSV_ASSIGNMENT_DELAY D_IN; end
             endcase
          end // else: !if(RST == `BSV_RESET_VALUE)
     end // always @ (posedge CLK)

   // Update the memory array  reset is OFF
   always @(posedge CLK `BSV_ARESET_EDGE_ARRAY)
     begin: array
`ifdef BSV_RESET_FIFO_ARRAY
        if (RST == `BSV_RESET_VALUE)
          begin: rst_array
             integer i;
             for (i = 0; i <= p2depth2 && p2depth > 2; i = i + 1)
               begin
                   arr[i]  <= `BSV_ASSIGNMENT_DELAY {p1width {1'b0}} ;
               end
          end // if (RST == `BSV_RESET_VALUE)
        else
`endif
         begin
            if (!CLR && ENQ && ((DEQ && !ring_empty) || (!DEQ && hasodata && not_ring_full)))
              begin
                 arr[tail] <= `BSV_ASSIGNMENT_DELAY D_IN;
              end
         end // else: !if(RST == `BSV_RESET_VALUE)
     end // always @ (posedge CLK)

   // synopsys translate_off
   always@(posedge CLK)
     begin: error_checks
        reg deqerror, enqerror ;

        deqerror =  0;
        enqerror = 0;
        if (RST == ! `BSV_RESET_VALUE)
           begin
              if ( ! EMPTY_N && DEQ )
                begin
                   deqerror = 1 ;
                   $display( "Warning: SizedFIFO: %m -- Dequeuing from empty fifo" ) ;
                end
              if ( ! FULL_N && ENQ && (!DEQ || guarded) )
                begin
                   enqerror =  1 ;
                   $display( "Warning: SizedFIFO: %m -- Enqueuing to a full fifo" ) ;
                end
           end
     end // block: error_checks
   // synopsys translate_on

   // synopsys translate_off
   // Some assertions about parameter values
   initial
     begin : parameter_assertions
        integer ok ;
        ok = 1 ;

        if ( p2depth <= 1)
          begin
             ok = 0;
             $display ( "Warning SizedFIFO: %m -- depth parameter increased from %0d to 2", p2depth);
          end

        if ( p3cntr_width <= 0 )
          begin
             ok = 0;
             $display ( "ERROR SizedFIFO: %m -- width parameter must be greater than 0" ) ;
          end

        if ( ok == 0 ) $finish ;

      end // initial begin
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


// A clock synchronization FIFO where the enqueue and dequeue sides are in
// different clock domains.
// The depth of the FIFO is strictly 1 element.   Implementation uses only
// 1 register to minimize hardware
// There are no restrictions w.r.t. clock frequencies
// FULL and EMPTY signal are pessimistic, that is, they are asserted
// immediately when the FIFO becomes FULL or EMPTY, but their deassertion
// is delayed due to synchronization latency.
module SyncFIFO1(
                 sCLK,
                 sRST,
                 dCLK,
                 sENQ,
                 sD_IN,
                 sFULL_N,
                 dDEQ,
                 dD_OUT,
                 dEMPTY_N
                 ) ;

   parameter                 dataWidth = 1 ;

   // input clock domain ports
   input                     sCLK ;
   input                     sRST ;
   input                     sENQ ;
   input [dataWidth -1 : 0]  sD_IN ;
   output                    sFULL_N ;

   // destination clock domain ports
   input                     dCLK ;
   input                     dDEQ ;
   output                    dEMPTY_N ;
   output [dataWidth -1 : 0] dD_OUT ;

   // FIFO DATA
   reg [dataWidth -1 : 0]    syncFIFO1Data ;

   // Reset generation
   wire                      dRST = sRST;

   // sCLK registers
   reg                       sEnqToggle,  sDeqToggle, sSyncReg1;
   // dCLK registers
   reg                       dEnqToggle,  dDeqToggle, dSyncReg1;

   // output assignment
   assign dD_OUT = syncFIFO1Data;
   assign dEMPTY_N = dEnqToggle != dDeqToggle;
   assign sFULL_N  = sEnqToggle == sDeqToggle;

   always @(posedge sCLK or `BSV_RESET_EDGE sRST) begin
      if (sRST == `BSV_RESET_VALUE) begin
         syncFIFO1Data <= `BSV_ASSIGNMENT_DELAY  {dataWidth {1'b0}};
         sEnqToggle    <= `BSV_ASSIGNMENT_DELAY  1'b0;
         sSyncReg1     <= `BSV_ASSIGNMENT_DELAY  1'b0;
         sDeqToggle    <= `BSV_ASSIGNMENT_DELAY  1'b1; // FIFO marked as full during reset
      end
      else begin
         if (sENQ && (sEnqToggle == sDeqToggle)) begin
            syncFIFO1Data <= `BSV_ASSIGNMENT_DELAY sD_IN;
            sEnqToggle    <= `BSV_ASSIGNMENT_DELAY ! sEnqToggle;
         end
         sSyncReg1  <= `BSV_ASSIGNMENT_DELAY dDeqToggle; // clock domain crossing
         sDeqToggle <= `BSV_ASSIGNMENT_DELAY sSyncReg1;
      end
   end

   always @(posedge dCLK or `BSV_RESET_EDGE dRST) begin
      if (dRST == `BSV_RESET_VALUE) begin
         dEnqToggle    <= `BSV_ASSIGNMENT_DELAY  1'b0;
         dSyncReg1     <= `BSV_ASSIGNMENT_DELAY  1'b0;
         dDeqToggle    <= `BSV_ASSIGNMENT_DELAY  1'b0;
      end
      else begin
         if (dDEQ && (dEnqToggle != dDeqToggle)) begin
            dDeqToggle    <= `BSV_ASSIGNMENT_DELAY ! dDeqToggle;
         end
         dSyncReg1  <= `BSV_ASSIGNMENT_DELAY sEnqToggle; // clock domain crossing
         dEnqToggle <= `BSV_ASSIGNMENT_DELAY dSyncReg1;
      end
   end

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin : initBlock
      syncFIFO1Data = {((dataWidth + 1)/2){2'b10}} ;
      sEnqToggle = 1'b0;
      sDeqToggle = 1'b0;
      sSyncReg1 = 1'b0;

      dEnqToggle = 1'b0;
      dDeqToggle = 1'b0;
      dSyncReg1 = 1'b0;
   end
   // synopsys translate_on
`endif // !`ifdef BSV_NO_INITIAL_BLOCKS

   // synopsys translate_off
   always@(posedge sCLK)
     begin: error_checks1
        reg enqerror ;
        enqerror = 0;
        if (sRST == ! `BSV_RESET_VALUE)
          begin
             if ( sENQ && (sEnqToggle != sDeqToggle)) begin
                enqerror = 1;
                $display( "Warning: SyncFIFO1: %m -- Enqueuing to a full fifo" ) ;
             end
          end
     end

   always@(posedge dCLK)
     begin: error_checks2
        reg deqerror ;
        deqerror = 0;
        if (dRST == ! `BSV_RESET_VALUE)
          begin
             if ( dDEQ && (dEnqToggle == dDeqToggle)) begin
                deqerror = 1;
                $display( "Warning: SyncFIFO1: %m -- Dequeuing from an empty full fifo" ) ;
             end
          end
     end // block: error_checks
   // synopsys translate_on

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_RESET_EDGE_HEAD or `BSV_RESET_EDGE dRST
`else
 `define BSV_RESET_EDGE_HEAD
`endif


// A clock synchronization FIFO where the enqueue and dequeue sides are in
// different clock domains.
// There are no restrictions w.r.t. clock frequencies
// The depth of the FIFO must be a power of 2 (2,4,8,...) since the
// indexing uses a Gray code counter.
// FULL and EMPTY signal are pessimistic, that is, they are asserted
// immediately when the FIFO becomes FULL or EMPTY, but their deassertion
// is delayed due to synchronization latency.
module SyncFIFO(
                sCLK,
                sRST,
                dCLK,
                sENQ,
                sD_IN,
                sFULL_N,
                dDEQ,
                dD_OUT,
                dEMPTY_N
                ) ;


   parameter                 dataWidth = 1 ;
   parameter                 depth = 2 ; // minimum 2
   parameter                 indxWidth = 1 ; // minimum 1

   // input clock domain ports
   input                     sCLK ;
   input                     sRST ;
   input                     sENQ ;
   input [dataWidth -1 : 0]  sD_IN ;
   output                    sFULL_N ;

   // destination clock domain ports
   input                     dCLK ;
   input                     dDEQ ;
   output                    dEMPTY_N ;
   output [dataWidth -1 : 0] dD_OUT ;

   // constants for bit masking of the gray code
   wire [indxWidth : 0]      msbset  = ~({(indxWidth + 1){1'b1}} >> 1) ;
   wire [indxWidth - 1 : 0]  msb2set = ~({(indxWidth + 0){1'b1}} >> 1) ;
   wire [indxWidth : 0]      msb12set = msbset | {1'b0, msb2set} ; // 'b11000...

   // FIFO Memory
   reg [dataWidth -1 : 0]    fifoMem [0: depth -1 ] ;
   reg [dataWidth -1 : 0]    dDoutReg ;

   // Enqueue Pointer support
   reg [indxWidth +1 : 0]    sGEnqPtr, sGEnqPtr1 ; // Flops
   reg                       sNotFullReg ;
   wire                      sNextNotFull, sFutureNotFull ;

   // Dequeue Pointer support
   reg [indxWidth+1 : 0]       dGDeqPtr, dGDeqPtr1 ; // Flops
   reg                       dNotEmptyReg ;
   wire                      dNextNotEmpty;

   // Reset generation
   wire                      dRST ;

   // flops to sychronize enqueue and dequeue point across domains
   reg [indxWidth : 0]       dSyncReg1, dEnqPtr ;
   reg [indxWidth : 0]       sSyncReg1, sDeqPtr ;

   wire [indxWidth - 1 :0]   sEnqPtrIndx, dDeqPtrIndx ;

   // Resets
   assign                    dRST = sRST ;

   // Outputs
   assign                    dD_OUT   = dDoutReg     ;
   assign                    dEMPTY_N = dNotEmptyReg ;
   assign                    sFULL_N  = sNotFullReg  ;

   // Indexes are truncated from the Gray counter with parity
   assign                    sEnqPtrIndx  = sGEnqPtr[indxWidth-1:0];
   assign                    dDeqPtrIndx  = dGDeqPtr[indxWidth-1:0];

   // Fifo memory write
   always @(posedge sCLK)
     begin
        if ( sENQ )
          fifoMem[sEnqPtrIndx] <= `BSV_ASSIGNMENT_DELAY sD_IN ;
     end // always @ (posedge sCLK)

   ////////////////////////////////////////////////////////////////////////
   // Enqueue Pointer and increment logic
   assign sNextNotFull   = (sGEnqPtr [indxWidth+1:1] ^ msb12set) != sDeqPtr ;
   assign sFutureNotFull = (sGEnqPtr1[indxWidth+1:1] ^ msb12set) != sDeqPtr ;

   always @(posedge sCLK or `BSV_RESET_EDGE sRST)
     begin
        if (sRST == `BSV_RESET_VALUE)
          begin
             sGEnqPtr    <= `BSV_ASSIGNMENT_DELAY {(indxWidth +2 ) {1'b0}} ;
             sGEnqPtr1   <= `BSV_ASSIGNMENT_DELAY { {indxWidth {1'b0}}, 2'b11} ;
             sNotFullReg <= `BSV_ASSIGNMENT_DELAY 1'b0 ; // Mark as full during reset to avoid spurious loads
          end // if (sRST == `BSV_RESET_VALUE)
        else
           begin
              if ( sENQ )
                begin
                   sGEnqPtr1   <= `BSV_ASSIGNMENT_DELAY incrGrayP( sGEnqPtr1 ) ;
                   sGEnqPtr    <= `BSV_ASSIGNMENT_DELAY sGEnqPtr1 ;
                   sNotFullReg <= `BSV_ASSIGNMENT_DELAY sFutureNotFull ;
                end // if ( sENQ )
              else
                begin
                   sNotFullReg <= `BSV_ASSIGNMENT_DELAY  sNextNotFull ;
                end // else: !if( sENQ )
           end // else: !if(sRST == `BSV_RESET_VALUE)
     end // always @ (posedge sCLK or `BSV_RESET_EDGE sRST)


   // Enqueue pointer synchronizer to dCLK
   always @(posedge dCLK  or `BSV_RESET_EDGE dRST)
     begin
        if (dRST == `BSV_RESET_VALUE)
          begin
             dSyncReg1 <= `BSV_ASSIGNMENT_DELAY {(indxWidth + 1) {1'b0}} ;
             dEnqPtr   <= `BSV_ASSIGNMENT_DELAY {(indxWidth + 1) {1'b0}} ;
          end // if (dRST == `BSV_RESET_VALUE)
        else
          begin
             dSyncReg1 <= `BSV_ASSIGNMENT_DELAY sGEnqPtr[indxWidth+1:1] ; // Clock domain crossing
             dEnqPtr   <= `BSV_ASSIGNMENT_DELAY dSyncReg1 ;
          end // else: !if(dRST == `BSV_RESET_VALUE)
     end // always @ (posedge dCLK  or `BSV_RESET_EDGE dRST)
   ////////////////////////////////////////////////////////////////////////


   ////////////////////////////////////////////////////////////////////////
   // Enqueue Pointer and increment logic
   assign dNextNotEmpty   = dGDeqPtr[indxWidth+1:1]  != dEnqPtr ;

   always @(posedge dCLK or `BSV_RESET_EDGE dRST)
     begin
        if (dRST == `BSV_RESET_VALUE)
          begin
             dGDeqPtr     <= `BSV_ASSIGNMENT_DELAY {(indxWidth + 2) {1'b0}} ;
             dGDeqPtr1    <= `BSV_ASSIGNMENT_DELAY {{indxWidth {1'b0}}, 2'b11 } ;
             dNotEmptyReg <= `BSV_ASSIGNMENT_DELAY 1'b0 ;
          end // if (dRST == `BSV_RESET_VALUE)
        else
           begin
              if ((!dNotEmptyReg || dDEQ) && dNextNotEmpty) begin
                 dGDeqPtr     <= `BSV_ASSIGNMENT_DELAY dGDeqPtr1 ;
                 dGDeqPtr1    <= `BSV_ASSIGNMENT_DELAY incrGrayP( dGDeqPtr1 );
                 dNotEmptyReg <= `BSV_ASSIGNMENT_DELAY 1'b1;
              end
              else if (dDEQ && !dNextNotEmpty) begin
                 dNotEmptyReg <= `BSV_ASSIGNMENT_DELAY 1'b0;
              end
           end // else: !if(dRST == `BSV_RESET_VALUE)
     end // always @ (posedge dCLK or `BSV_RESET_EDGE dRST)


   always @(posedge dCLK `BSV_RESET_EDGE_HEAD)
     begin
`ifdef  BSV_RESET_FIFO_HEAD
        if (dRST == `BSV_RESET_VALUE)
          begin
             dDoutReg    <= `BSV_ASSIGNMENT_DELAY {dataWidth {1'b0}} ;
          end // if (dRST == `BSV_RESET_VALUE)
        else
`endif
          begin
             if ((!dNotEmptyReg || dDEQ) && dNextNotEmpty) begin
                dDoutReg     <= `BSV_ASSIGNMENT_DELAY fifoMem[dDeqPtrIndx] ;
             end
          end
     end

    // Dequeue pointer synchronized to sCLK
    always @(posedge sCLK  or `BSV_RESET_EDGE sRST)
      begin
         if (sRST == `BSV_RESET_VALUE)
           begin
              sSyncReg1 <= `BSV_ASSIGNMENT_DELAY {(indxWidth + 1) {1'b0}} ;
              sDeqPtr   <= `BSV_ASSIGNMENT_DELAY {(indxWidth + 1) {1'b0}} ; // When reset mark as not empty
           end // if (sRST == `BSV_RESET_VALUE)
         else
           begin
              sSyncReg1 <= `BSV_ASSIGNMENT_DELAY dGDeqPtr[indxWidth+1:1] ; // clock domain crossing
              sDeqPtr   <= `BSV_ASSIGNMENT_DELAY sSyncReg1 ;
           end // else: !if(sRST == `BSV_RESET_VALUE)
      end // always @ (posedge sCLK  or `BSV_RESET_EDGE sRST)
   ////////////////////////////////////////////////////////////////////////

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin : initBlock
        integer i ;

        // initialize the FIFO memory with aa's
        for (i = 0; i < depth; i = i + 1)
          begin
             fifoMem[i] = {((dataWidth + 1)/2){2'b10}} ;
          end
        dDoutReg     = {((dataWidth + 1)/2){2'b10}} ;

        // initialize the pointer
        sGEnqPtr = {((indxWidth + 2)/2){2'b10}} ;
        sGEnqPtr1 = sGEnqPtr ;
        sNotFullReg = 1'b0 ;

        dGDeqPtr = sGEnqPtr ;
        dGDeqPtr1 = sGEnqPtr ;
        dNotEmptyReg = 1'b0;


        // initialize other registers
        sSyncReg1 = sGEnqPtr ;
        sDeqPtr   = sGEnqPtr ;
        dSyncReg1 = sGEnqPtr ;
        dEnqPtr   = sGEnqPtr ;
     end // block: initBlock
   // synopsys translate_on



   // synopsys translate_off
   initial
     begin : parameter_assertions
        integer ok ;
        integer i, expDepth ;

        ok = 1;
        expDepth = 1 ;

        // calculate x = 2 ** (indxWidth - 1)
        for( i = 0 ; i < indxWidth ; i = i + 1 )
          begin
             expDepth = expDepth * 2 ;
          end // for ( i = 0 ; i < indxWidth ; i = i + 1 )

        if ( expDepth != depth )
          begin
             ok = 0;
             $display ( "ERROR SyncFiFO.v: index size and depth do not match;" ) ;
             $display ( "\tdepth must equal 2 ** index size. expected %0d", expDepth );
          end

        #0
        if ( ok == 0 ) $finish ;

      end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

   function [indxWidth+1:0] incrGrayP ;
      input [indxWidth+1:0] grayPin;

      begin: incrGrayPBlock
         reg [indxWidth :0] g;
         reg                p ;
         reg [indxWidth :0] i;

         g = grayPin[indxWidth+1:1];
         p = grayPin[0];
         i = incrGray (g,p);
         incrGrayP = {i,~p};
      end
   endfunction
   function [indxWidth:0] incrGray ;
      input [indxWidth:0] grayin;
      input parity ;

      begin: incrGrayBlock
         integer               i;
         reg [indxWidth: 0]    tempshift;
         reg [indxWidth: 0]    flips;

         flips[0] = ! parity ;
         for ( i = 1 ; i < indxWidth ; i = i+1 )
           begin
              tempshift = grayin << (2 + indxWidth - i ) ;
              flips[i]  = parity & grayin[i-1] & ~(| tempshift ) ;
           end
         tempshift = grayin << 2 ;
         flips[indxWidth] = parity & ~(| tempshift ) ;

         incrGray = flips ^ grayin ;
      end
   endfunction

endmodule // FIFOSync


`ifdef testBluespec
module testSyncFIFO() ;
   parameter dsize = 8;
   parameter fifodepth = 32;
   parameter fifoidx = 5;

   wire      sCLK,  dCLK, dRST ;
   wire      sENQ, dDEQ;
   wire      sFULL_N, dEMPTY_N ;
   wire [dsize -1:0] sDIN, dDOUT ;

   reg [dsize -1:0]  sCNT, dCNT ;
   reg sRST, sCLR ;

   ClockGen#(15,14,10)  sc( sCLK );
   ClockGen#(11,12,2600)  dc( dCLK );

   initial
     begin
        sCNT = 0;
        dCNT = 0;
        sCLR = 1'b0 ;

        sRST = `BSV_RESET_VALUE ;
        $display( "running test" ) ;

        $dumpfile("SyncFIFO.vcd");
        $dumpvars(5,testSyncFIFO) ;
        $dumpon ;
        #200 ;
        sRST = !`BSV_RESET_VALUE ;


        #100000 $finish ;
     end // initial begin
   initial
     begin
        #50000 ;
        @(posedge sCLK ) ;
        sCLR <= `BSV_ASSIGNMENT_DELAY 1'b1 ;
        @(posedge sCLK ) ;
        sCLR <= `BSV_ASSIGNMENT_DELAY 1'b0 ;

      end

   SyncFIFO #(dsize,fifodepth,fifoidx)
     dut( sCLK, sRST, dCLK, sENQ, sDIN,
          sFULL_N, // sCLR,
          dDEQ, dDOUT, dEMPTY_N );

   assign sDIN = sCNT ;
   assign sENQ = sFULL_N ;


   always @(posedge sCLK)
     begin
        if (sENQ )
          begin
             sCNT <= `BSV_ASSIGNMENT_DELAY sCNT + 1;
          end
      end // always @ (posedge sCLK)

   assign dDEQ = dEMPTY_N ;

   always @(posedge dCLK)
     begin
        if (dDEQ )
           begin
              $display( "dequeing %d", dDOUT ) ;
           end
     end // always @ (posedge dCLK)

endmodule // testSyncFIFO
`endif
// Copyright (c) 2000-2013 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


//
// Transfer takes 2 dCLK to see data,
// sRDY recovers takes 2 dCLK + 2 sCLK
module SyncHandshake(
                     sCLK,
                     sRST,
                     dCLK,
                     sEN,
                     sRDY,
                     dPulse
                     );
   parameter init = 1'b0;
   parameter delayreturn = 1'b0;

   // Source clock port signal
   input     sCLK ;
   input     sRST ;
   input     sEN ;
   output    sRDY ;

   // Destination clock port signal
   input     dCLK ;
   output    dPulse ;

   // Flops to hold data
   reg       dSyncReg1, dSyncReg2 ;
   reg       dLastState ;
   reg       sToggleReg ;
   reg       sSyncReg1, sSyncReg2 ;

   // Output signal
   assign    dPulse = dSyncReg2 != dLastState ;
   assign    sRDY = sSyncReg2 == sToggleReg;
   wire      ackValue = delayreturn ? dLastState : dSyncReg2 ;

   always @(posedge sCLK or `BSV_RESET_EDGE sRST)
     begin
        if (sRST == `BSV_RESET_VALUE)
           begin
              sSyncReg1  <= `BSV_ASSIGNMENT_DELAY ! init ; // Reset hi so sRDY is low during reset
              sSyncReg2  <= `BSV_ASSIGNMENT_DELAY ! init ;
              sToggleReg <= `BSV_ASSIGNMENT_DELAY init ;
           end
        else
           begin

              // hadshake return synchronizer
              sSyncReg1 <= `BSV_ASSIGNMENT_DELAY ackValue ;// clock domain crossing
              sSyncReg2 <= `BSV_ASSIGNMENT_DELAY sSyncReg1 ;

              // Pulse send
              if ( sEN )
                begin
                   sToggleReg <= `BSV_ASSIGNMENT_DELAY ! sToggleReg ;
                end // if ( sEN )

           end
     end // always @ (posedge sCLK or `BSV_RESET_EDGE sRST)

   always @(posedge dCLK or `BSV_RESET_EDGE sRST)
     begin
        if (sRST == `BSV_RESET_VALUE)
          begin
             dSyncReg1  <= `BSV_ASSIGNMENT_DELAY init;
             dSyncReg2  <= `BSV_ASSIGNMENT_DELAY init;
             dLastState <= `BSV_ASSIGNMENT_DELAY init ;
          end
        else
           begin
              dSyncReg1 <= `BSV_ASSIGNMENT_DELAY sToggleReg ;// domain crossing
              dSyncReg2 <= `BSV_ASSIGNMENT_DELAY dSyncReg1 ;
              dLastState <= `BSV_ASSIGNMENT_DELAY dSyncReg2 ;
           end
     end // always @ (posedge dCLK or `BSV_RESET_EDGE sRST)

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
      begin
         dSyncReg1 = init ;
         dSyncReg2 = init ;
         dLastState = init ;

         sToggleReg = init ;
         sSyncReg1 = ! init ;
         sSyncReg2 = ! init ;

      end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule // HandshakeSync

// Copyright (c) 2000-2013 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif


// A register synchronization module across clock domains.
// Uses a Handshake Pulse protocol to trigger the load on
// destination side registers
// Transfer takes 3 dCLK for destination side to see data,
// sRDY recovers takes 3 dCLK + 3 sCLK
module SyncRegister(
                    sCLK,
                    sRST,
                    dCLK,
                    sEN,
                    sRDY,
                    sD_IN,
                    dD_OUT
                    );
   parameter             width = 1 ;
   parameter             init = { width {1'b0 }} ;

   // Source clock domain ports
   input                 sCLK ;
   input                 sRST ;
   input                 sEN ;
   input [width -1 : 0]  sD_IN ;
   output                sRDY ;

   // Destination clock domain ports
   input                 dCLK ;
   output [width -1 : 0] dD_OUT ;

   wire                  dPulse ;
   reg [width -1 : 0]    sDataSyncIn ;
   reg [width -1 : 0]    dD_OUT ;

   // instantiate a Handshake Sync
   SyncHandshake #(.init(0),.delayreturn(1))
   sync( .sCLK(sCLK), .sRST(sRST),
         .dCLK(dCLK),
         .sEN(sEN), .sRDY(sRDY),
         .dPulse(dPulse) ) ;

   always @(posedge sCLK or `BSV_RESET_EDGE sRST)
      begin
         if (sRST == `BSV_RESET_VALUE)
           begin
              sDataSyncIn <= `BSV_ASSIGNMENT_DELAY init ;
           end // if (sRST == `BSV_RESET_VALUE)
         else
           begin
              if ( sEN )
                begin
                   sDataSyncIn <= `BSV_ASSIGNMENT_DELAY sD_IN ;
                end // if ( sEN )
           end // else: !if(sRST == `BSV_RESET_VALUE)
      end // always @ (posedge sCLK or `BSV_RESET_EDGE sRST)


   // Transfer the data to destination domain when dPulsed is asserted.
   // Setup and hold time are assured since at least 2 dClks occured since
   // sDataSyncIn have been written.
   always @(posedge dCLK or `BSV_RESET_EDGE sRST)
      begin
         if (sRST == `BSV_RESET_VALUE)
           begin
              dD_OUT <= `BSV_ASSIGNMENT_DELAY init ;
           end // if (sRST == `BSV_RESET_VALUE)
         else
            begin
               if ( dPulse )
                 begin
                    dD_OUT <= `BSV_ASSIGNMENT_DELAY sDataSyncIn ;// clock domain crossing
                 end // if ( dPulse )
            end // else: !if(sRST == `BSV_RESET_VALUE)
      end // always @ (posedge dCLK or `BSV_RESET_EDGE sRST)


`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
      begin
         sDataSyncIn = {((width + 1)/2){2'b10}} ;
         dD_OUT      = {((width + 1)/2){2'b10}} ;
      end // initial begin
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS


endmodule // RegisterSync



`ifdef testBluespec
module testSyncRegister() ;
   parameter dsize = 8;

   wire      sCLK, sRST, dCLK ;
   wire      sEN ;
   wire      sRDY ;

   reg [dsize -1:0]  sCNT ;
   wire [dsize -1:0] sDIN, dDOUT ;

   ClockGen#(20,9,10)  sc( sCLK );
   ClockGen#(11,12,26)  dc( dCLK );

   initial
     begin
        sCNT = 0;

        $dumpfile("SyncRegister.dump");
        $dumpvars(5) ;
        $dumpon ;
        #100000 $finish ;
     end

   SyncRegister #(dsize)
     dut( sCLK, sRST, dCLK,
          sEN, sRDY, sDIN,
          dDOUT ) ;


   assign sDIN = sCNT ;
   assign sEN = sRDY ;

   always @(posedge sCLK)
     begin
        if (sRDY )
          begin
             sCNT <= `BSV_ASSIGNMENT_DELAY sCNT + 1;
          end
      end // always @ (posedge sCLK)



endmodule // testSyncFIFO
`endif



// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif



module SyncReset0 (
		   IN_RST,
		   OUT_RST
		   );

   input   IN_RST ;
   output  OUT_RST ;

   assign  OUT_RST = IN_RST ;

endmodule

// Copyright (c) 2000-2012 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif



// A synchronization module for resets.   Output resets are held for
// RSTDELAY+1 cycles, RSTDELAY >= 0.  Reset assertion is asynchronous,
// while deassertion is synchronized to the clock.
module SyncResetA (
                   IN_RST,
                   CLK,
                   OUT_RST
                   );

   parameter          RSTDELAY = 1  ; // Width of reset shift reg

   input              CLK ;
   input              IN_RST ;
   output             OUT_RST ;

   reg [RSTDELAY:0]   reset_hold ;
   wire [RSTDELAY+1:0] next_reset = {reset_hold, ~ `BSV_RESET_VALUE} ;

   assign  OUT_RST = reset_hold[RSTDELAY] ;

   always @( posedge CLK or `BSV_RESET_EDGE IN_RST )
     begin
        if (IN_RST == `BSV_RESET_VALUE)
           begin
              reset_hold <= `BSV_ASSIGNMENT_DELAY {RSTDELAY+1 {`BSV_RESET_VALUE}} ;
           end
        else
          begin
             reset_hold <= `BSV_ASSIGNMENT_DELAY next_reset[RSTDELAY:0];
          end
     end // always @ ( posedge CLK or  `BSV_RESET_EDGE IN_RST )

`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
     begin
        #0 ;
        // initialize out of reset forcing the designer to do one
        reset_hold = {(RSTDELAY + 1) {~ `BSV_RESET_VALUE}} ;
     end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule // SyncResetA

// Copyright (c) 2000-2009 Bluespec, Inc.

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
// $Revision$
// $Date$

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif

// A separate module which instantiates a simple clock muxing primitive.
// The primitive includes an internal register which maintains the selector
// state.
module UngatedClockMux(
                CLK,
                SELECT,
                SELECT_ENABLE,
                A_CLK,
                B_CLK,
                CLK_OUT
               ) ;

   input            CLK;
   input            SELECT;
   input            SELECT_ENABLE;

   input            A_CLK;
   input            B_CLK;

   output           CLK_OUT;

   reg sel_reg;

   assign CLK_OUT = sel_reg == 1'b1 ? A_CLK : B_CLK ;
   

   always @(posedge CLK)
   begin
     if (SELECT_ENABLE)
       sel_reg <= SELECT;
   end

      
`ifdef BSV_NO_INITIAL_BLOCKS
`else // not BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial
      begin
         #0 ;
         sel_reg  = 1'b0 ;
      end
   // synopsys translate_on
`endif // BSV_NO_INITIAL_BLOCKS

endmodule                
